
-- ARCHIVO AUTOGENERADO CON model/tensorflow_model.py

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.perceptron_package.perceptron_input;

package mnist_inputs_7 is
    function GetInputs(Dummy: natural)
    return perceptron_input;
end package mnist_inputs_7;

package body mnist_inputs_7 is
    function GetInputs(Dummy: natural) return perceptron_input is
        variable pesos_i : perceptron_input(63 downto 0);
    begin
	pesos_i(0) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(1) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(2) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(3) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(4) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(5) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(6) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(7) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(8) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(9) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(10) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(11) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(12) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(13) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(14) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(15) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(16) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(17) := b"0000000000000000_0000000000000001_0000000000000000_0000000000000000"; -- 1.0
	pesos_i(18) := b"0000000000000000_0000000000000000_1111111101000111_1100011100111100"; -- 0.997188999300896
	pesos_i(19) := b"0000000000000000_0000000000000000_1000110100001010_0011010011111110"; -- 0.5509369964982768
	pesos_i(20) := b"0000000000000000_0000000000000000_1001011110011000_1110000101010000"; -- 0.5921765155566483
	pesos_i(21) := b"0000000000000000_0000000000000000_1010000011001010_1110100100000111"; -- 0.6280961648762619
	pesos_i(22) := b"0000000000000000_0000000000000000_1111010100110100_0001101001111010"; -- 0.9578262852211513
	pesos_i(23) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(24) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(25) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(26) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(27) := b"0000000000000000_0000000000000000_0000010000100101_1111001010000000"; -- 0.016204029308772846
	pesos_i(28) := b"0000000000000000_0000000000000000_0001000110010011_1001010010001111"; -- 0.0686581467312056
	pesos_i(29) := b"0000000000000000_0000000000000000_1011001001001011_0011101000011110"; -- 0.6964603732981679
	pesos_i(30) := b"0000000000000000_0000000000000000_0100100110001111_1010000110001011"; -- 0.2873478855663454
	pesos_i(31) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(32) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(33) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(34) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(35) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(36) := b"0000000000000000_0000000000000000_0101101100101101_1001001010100101"; -- 0.35616413616812903
	pesos_i(37) := b"0000000000000000_0000000000000000_0101100010011001_1001101010000110"; -- 0.3460938051358994
	pesos_i(38) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(39) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(40) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(41) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(42) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(43) := b"0000000000000000_0000000000000000_0001001010101010_1100001101000000"; -- 0.07291813188947781
	pesos_i(44) := b"0000000000000000_0000000000000000_1011000111110110_0100000000100110"; -- 0.6951637356534567
	pesos_i(45) := b"0000000000000000_0000000000000000_0000011010010000_0001111001101001"; -- 0.02563657815821477
	pesos_i(46) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(47) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(48) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(49) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(50) := b"0000000000000000_0000000000000000_0000000110111100_1001000111100110"; -- 0.006783598634699972
	pesos_i(51) := b"0000000000000000_0000000000000000_1001101110001111_0000010110111110"; -- 0.6076510990789817
	pesos_i(52) := b"0000000000000000_0000000000000000_0010111100111100_1001111101000000"; -- 0.18451876934011505
	pesos_i(53) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(54) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(55) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(56) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(57) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(58) := b"0000000000000000_0000000000000000_0001001100011010_0100010011100101"; -- 0.0746195849816997
	pesos_i(59) := b"0000000000000000_0000000000000000_1001000100110000_0010011101111110"; -- 0.5671410258070496
	pesos_i(60) := b"0000000000000000_0000000000000000_0000010101111110_0001111001101101"; -- 0.021455670853501748
	pesos_i(61) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(62) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(63) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0

    return pesos_i;
    end function;
end package body mnist_inputs_7;
    