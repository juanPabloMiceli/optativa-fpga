
-- ARCHIVO AUTOGENERADO CON model/tensorflow_model.py

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.perceptron_package.perceptron_input;

package mnist_inputs_5 is
    function GetInputs(Dummy: natural)
    return perceptron_input;
end package mnist_inputs_5;

package body mnist_inputs_5 is
    function GetInputs(Dummy: natural) return perceptron_input is
        variable pesos_i : perceptron_input(63 downto 0);
    begin
	pesos_i(0) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(1) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(2) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(3) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(4) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(5) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(6) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(7) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(8) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(9) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(10) := b"0000000000000000_0000000000000000_0000101001100100_1101011000001010"; -- 0.04060113651690523
	pesos_i(11) := b"0000000000000000_0000000000000000_0010100100110001_1111101100000111"; -- 0.1609188931140404
	pesos_i(12) := b"0000000000000000_0000000000000000_0100111010111010_0111001011101000"; -- 0.30753248381292
	pesos_i(13) := b"0000000000000000_0000000000000000_0111110000001100_0011001010100011"; -- 0.4845611236320715
	pesos_i(14) := b"0000000000000000_0000000000000000_1111111100001001_1001111110001001"; -- 0.996240588195683
	pesos_i(15) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(16) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(17) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(18) := b"0000000000000000_0000000000000000_1001010011111010_1010011010001000"; -- 0.5819496234089749
	pesos_i(19) := b"0000000000000000_0000000000000000_1011000001110000_1010001001000001"; -- 0.6892186554129655
	pesos_i(20) := b"0000000000000000_0000000000000000_0111110010010100_1100000100010110"; -- 0.48664480955011513
	pesos_i(21) := b"0000000000000000_0000000000000000_0011101011100100_0010110010111010"; -- 0.23004416980512485
	pesos_i(22) := b"0000000000000000_0000000000000000_0001011000101101_0101101111001001"; -- 0.086629616364842
	pesos_i(23) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(24) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(25) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(26) := b"0000000000000000_0000000000000000_0000000100100111_1010011000000001"; -- 0.004511237390767247
	pesos_i(27) := b"0000000000000000_0000000000000000_0110001010110110_1000111010100111"; -- 0.3855981023676062
	pesos_i(28) := b"0000000000000000_0000000000000000_0010011111001011_1111011010010010"; -- 0.155455980828509
	pesos_i(29) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(30) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(31) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(32) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(33) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(34) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(35) := b"0000000000000000_0000000000000000_0000010101110000_1101110110001000"; -- 0.021253438713175147
	pesos_i(36) := b"0000000000000000_0000000000000000_0111100100011110_1101100000101011"; -- 0.47312689817372305
	pesos_i(37) := b"0000000000000000_0000000000000000_1000010011010001_1001010111100101"; -- 0.518823021262622
	pesos_i(38) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(39) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(40) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(41) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(42) := b"0000000000000000_0000000000000000_0000000100100111_1010011000000001"; -- 0.004511237390767247
	pesos_i(43) := b"0000000000000000_0000000000000000_0011000110111110_1100010011011101"; -- 0.19431715394902993
	pesos_i(44) := b"0000000000000000_0000000000000000_1010000000001101_0101010010000001"; -- 0.625203401158134
	pesos_i(45) := b"0000000000000000_0000000000000000_1010101001101000_1010110011111111"; -- 0.6656597253935528
	pesos_i(46) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(47) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(48) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(49) := b"0000000000000000_0000000000000000_1110110110110000_1010010111111110"; -- 0.9284766908852593
	pesos_i(50) := b"0000000000000000_0000000000000000_1100110110010001_0110110010111100"; -- 0.8030002555565701
	pesos_i(51) := b"0000000000000000_0000000000000000_1000111100000100_0111010111111100"; -- 0.558661817603461
	pesos_i(52) := b"0000000000000000_0000000000000000_0010110000011111_0101100110111000"; -- 0.17235337004899912
	pesos_i(53) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(54) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(55) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(56) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(57) := b"0000000000000000_0000000000000000_0101111100010011_0111010110011001"; -- 0.3713906763541037
	pesos_i(58) := b"0000000000000000_0000000000000000_0001111100101110_1000001000011101"; -- 0.12180340955071568
	pesos_i(59) := b"0000000000000000_0000000000000000_0000001001010100_1111000100111010"; -- 0.009108616591360778
	pesos_i(60) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(61) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(62) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(63) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0

    return pesos_i;
    end function;
end package body mnist_inputs_5;
    