
-- ARCHIVO AUTOGENERADO CON model/tensorflow_model.py

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.perceptron_package.perceptron_input;

package mnist_weights is
    function GetWeights(Dummy: natural)
    return perceptron_input;
end package mnist_weights;

package body mnist_weights is
    function GetWeights(Dummy: natural) return perceptron_input is
        variable pesos_i : perceptron_input(9471 downto 0);
    begin
	pesos_i(0) := b"1111111111111111_1111111111111111_1101010001010001_0010100111000000"; -- -0.17063654959201813
	pesos_i(1) := b"1111111111111111_1111111111111111_1111101100011001_0010111100000000"; -- -0.019146978855133057
	pesos_i(2) := b"1111111111111111_1111111111111111_1111111111010001_1011000110011110"; -- -0.0007065762765705585
	pesos_i(3) := b"0000000000000000_0000000000000000_0000011000100101_0101100010010000"; -- 0.02400735393166542
	pesos_i(4) := b"1111111111111111_1111111111111111_1101111110010000_1001111110000000"; -- -0.12669947743415833
	pesos_i(5) := b"1111111111111111_1111111111111111_1110011000111100_1000100101000000"; -- -0.10063879191875458
	pesos_i(6) := b"0000000000000000_0000000000000000_0001011111010010_1110101000100000"; -- 0.09306205064058304
	pesos_i(7) := b"0000000000000000_0000000000000000_0001100111111100_1101110111100000"; -- 0.10151468962430954
	pesos_i(8) := b"1111111111111111_1111111111111111_1101001111111111_1001000001000000"; -- -0.17188166081905365
	pesos_i(9) := b"0000000000000000_0000000000000000_0010010011011001_0100110110000000"; -- 0.1439407765865326
	pesos_i(10) := b"0000000000000000_0000000000000000_0001001011111100_1101110110000000"; -- 0.07417091727256775
	pesos_i(11) := b"1111111111111111_1111111111111111_1101101101101100_0001000111000000"; -- -0.14288224279880524
	pesos_i(12) := b"0000000000000000_0000000000000000_0100000110111001_0111111000000000"; -- 0.2567366361618042
	pesos_i(13) := b"0000000000000000_0000000000000000_0011101001011100_1000110011000000"; -- 0.22797469794750214
	pesos_i(14) := b"0000000000000000_0000000000000000_0011111011111100_0000111101000000"; -- 0.24603362381458282
	pesos_i(15) := b"1111111111111111_1111111111111111_1110101111000101_1010110111000000"; -- -0.07901491224765778
	pesos_i(16) := b"1111111111111111_1111111111111111_1011110001001001_1100100110000000"; -- -0.26449909806251526
	pesos_i(17) := b"0000000000000000_0000000000000000_0000101001001010_0110110001010000"; -- 0.040198106318712234
	pesos_i(18) := b"1111111111111111_1111111111111111_1111100101101110_1001001100111000"; -- -0.025656508281826973
	pesos_i(19) := b"0000000000000000_0000000000000000_0001100010101100_1010100100100000"; -- 0.09638459235429764
	pesos_i(20) := b"0000000000000000_0000000000000000_0001100110010101_1000111100100000"; -- 0.09993834048509598
	pesos_i(21) := b"1111111111111111_1111111111111111_1101111101011100_1101000110000000"; -- -0.12748995423316956
	pesos_i(22) := b"1111111111111111_1111111111111111_1110110000000011_0011101000000000"; -- -0.07807576656341553
	pesos_i(23) := b"1111111111111111_1111111111111111_1110110001000001_0011101100100000"; -- -0.07712965458631516
	pesos_i(24) := b"1111111111111111_1111111111111111_1100111010101011_1010001110000000"; -- -0.19269350171089172
	pesos_i(25) := b"1111111111111111_1111111111111111_1111010100110111_1000111000000000"; -- -0.042121052742004395
	pesos_i(26) := b"1111111111111111_1111111111111111_1111100001101101_0110011000001000"; -- -0.02958071045577526
	pesos_i(27) := b"0000000000000000_0000000000000000_0010001101000110_0111110010000000"; -- 0.13779428601264954
	pesos_i(28) := b"0000000000000000_0000000000000000_0010011111010010_0101010001000000"; -- 0.15555311739444733
	pesos_i(29) := b"1111111111111111_1111111111111111_1110101000011001_1000000001000000"; -- -0.08554838597774506
	pesos_i(30) := b"0000000000000000_0000000000000000_0001010100110100_0110111000000000"; -- 0.08283126354217529
	pesos_i(31) := b"0000000000000000_0000000000000000_0001011011100110_0011010001100000"; -- 0.08945014327764511
	pesos_i(32) := b"1111111111111111_1111111111111111_1110011100100011_1000110011100000"; -- -0.09711379557847977
	pesos_i(33) := b"0000000000000000_0000000000000000_0010110000100000_1101010000000000"; -- 0.17237591743469238
	pesos_i(34) := b"1111111111111111_1111111111111111_1111111000000101_1110000111001100"; -- -0.007722747512161732
	pesos_i(35) := b"0000000000000000_0000000000000000_0000011110011101_1000010111001000"; -- 0.029747353866696358
	pesos_i(36) := b"1111111111111111_1111111111111111_1111001001110110_1010100111010000"; -- -0.05287684127688408
	pesos_i(37) := b"0000000000000000_0000000000000000_0000000011110100_1100111001111000"; -- 0.003735451027750969
	pesos_i(38) := b"1111111111111111_1111111111111111_1110000011100000_1100100010100000"; -- -0.12157007306814194
	pesos_i(39) := b"0000000000000000_0000000000000000_0001100110000110_0011110011000000"; -- 0.0997045487165451
	pesos_i(40) := b"0000000000000000_0000000000000000_0001000100010001_0000011000000000"; -- 0.06666600704193115
	pesos_i(41) := b"0000000000000000_0000000000000000_0001011010000101_0011011010000000"; -- 0.08797016739845276
	pesos_i(42) := b"0000000000000000_0000000000000000_0001111000110111_0000001001000000"; -- 0.11802686750888824
	pesos_i(43) := b"0000000000000000_0000000000000000_0001101110100010_0010000111100000"; -- 0.10794269293546677
	pesos_i(44) := b"0000000000000000_0000000000000000_0001100111110111_0101011101000000"; -- 0.10143037140369415
	pesos_i(45) := b"0000000000000000_0000000000000000_0010000011110101_1110101111000000"; -- 0.1287524551153183
	pesos_i(46) := b"0000000000000000_0000000000000000_0001001001000101_1011010101000000"; -- 0.07137615978717804
	pesos_i(47) := b"1111111111111111_1111111111111111_1111100010001110_1101100110001000"; -- -0.029070286080241203
	pesos_i(48) := b"0000000000000000_0000000000000000_0100100010111000_1010011000000000"; -- 0.2840675115585327
	pesos_i(49) := b"1111111111111111_1111111111111111_1111101000010111_1010000101101000"; -- -0.023076927289366722
	pesos_i(50) := b"1111111111111111_1111111111111111_1111101110101010_0001010100111000"; -- -0.016935991123318672
	pesos_i(51) := b"0000000000000000_0000000000000000_0011001000010100_0110100010000000"; -- 0.19562390446662903
	pesos_i(52) := b"0000000000000000_0000000000000000_0010011000011100_0100111001000000"; -- 0.14886941015720367
	pesos_i(53) := b"0000000000000000_0000000000000000_0000111110110111_1111100110000000"; -- 0.06140097975730896
	pesos_i(54) := b"1111111111111111_1111111111111111_1110010001111011_1100010101000000"; -- -0.10748641192913055
	pesos_i(55) := b"0000000000000000_0000000000000000_0000110010110110_0010100111000000"; -- 0.04965458810329437
	pesos_i(56) := b"0000000000000000_0000000000000000_0001011111111001_1100110111000000"; -- 0.09365545213222504
	pesos_i(57) := b"0000000000000000_0000000000000000_0000111111000100_1110110000000000"; -- 0.06159853935241699
	pesos_i(58) := b"0000000000000000_0000000000000000_0001011010100110_0100001100000000"; -- 0.08847445249557495
	pesos_i(59) := b"0000000000000000_0000000000000000_0000000111011001_0000111101101110"; -- 0.007218326907604933
	pesos_i(60) := b"1111111111111111_1111111111111111_1111100010111111_0100111100010000"; -- -0.028330858796834946
	pesos_i(61) := b"0000000000000000_0000000000000000_0010011011010001_0101111000000000"; -- 0.1516321897506714
	pesos_i(62) := b"1111111111111111_1111111111111111_1100000001000000_0101100011000000"; -- -0.24901814758777618
	pesos_i(63) := b"1111111111111111_1111111111111111_1110110011100010_1001101101000000"; -- -0.07466726005077362
	pesos_i(64) := b"1111111111111111_1111111111111111_1111111010011110_1001011110000010"; -- -0.005392580758780241
	pesos_i(65) := b"0000000000000000_0000000000000000_0001000011011001_1001011001100000"; -- 0.0658201202750206
	pesos_i(66) := b"0000000000000000_0000000000000000_0011110111110010_1101001001000000"; -- 0.24198640882968903
	pesos_i(67) := b"1111111111111111_1111111111111111_1101101100010100_0000101010000000"; -- -0.14422544836997986
	pesos_i(68) := b"1111111111111111_1111111111111111_1111001111011011_0111001111000000"; -- -0.04743267595767975
	pesos_i(69) := b"0000000000000000_0000000000000000_0000111000011010_0000000001110000"; -- 0.05508425459265709
	pesos_i(70) := b"0000000000000000_0000000000000000_0001101111100010_1101001111000000"; -- 0.10892985761165619
	pesos_i(71) := b"1111111111111111_1111111111111111_1111001000101111_1101000010000000"; -- -0.05395790934562683
	pesos_i(72) := b"0000000000000000_0000000000000000_0011001001010101_0010101011000000"; -- 0.19661204516887665
	pesos_i(73) := b"0000000000000000_0000000000000000_0011001001011011_1111011101000000"; -- 0.19671578705310822
	pesos_i(74) := b"0000000000000000_0000000000000000_0001011110100000_1011000100000000"; -- 0.09229570627212524
	pesos_i(75) := b"0000000000000000_0000000000000000_0001110000110000_0010010001000000"; -- 0.11010958254337311
	pesos_i(76) := b"0000000000000000_0000000000000000_0011011101110100_0011010111000000"; -- 0.21661697328090668
	pesos_i(77) := b"1111111111111111_1111111111111111_1100100001001100_1010111011000000"; -- -0.2175799161195755
	pesos_i(78) := b"0000000000000000_0000000000000000_0000000110011010_0001000010100010"; -- 0.006257094908505678
	pesos_i(79) := b"0000000000000000_0000000000000000_0010010010001100_0101101111000000"; -- 0.14276669919490814
	pesos_i(80) := b"1111111111111111_1111111111111111_1110110111010110_0101001011000000"; -- -0.07094843685626984
	pesos_i(81) := b"0000000000000000_0000000000000000_0100000011110001_1000010000000000"; -- 0.25368523597717285
	pesos_i(82) := b"1111111111111111_1111111111111111_1111010100101001_1000001011100000"; -- -0.04233533889055252
	pesos_i(83) := b"0000000000000000_0000000000000000_0011011010010101_0101010000000000"; -- 0.21321606636047363
	pesos_i(84) := b"0000000000000000_0000000000000000_0000100001011000_1100010011100000"; -- 0.032604508101940155
	pesos_i(85) := b"1111111111111111_1111111111111111_1110110101111011_0010010000100000"; -- -0.07233976572751999
	pesos_i(86) := b"0000000000000000_0000000000000000_0001000000000011_1110110000100000"; -- 0.06255985051393509
	pesos_i(87) := b"1111111111111111_1111111111111111_1111110000111001_1110000111101000"; -- -0.01474178396165371
	pesos_i(88) := b"0000000000000000_0000000000000000_0011010001110010_1011111001000000"; -- 0.20487584173679352
	pesos_i(89) := b"0000000000000000_0000000000000000_0000010011000001_0001010011101000"; -- 0.018571192398667336
	pesos_i(90) := b"1111111111111111_1111111111111111_1101101110101110_0010010111000000"; -- -0.14187397062778473
	pesos_i(91) := b"1111111111111111_1111111111111111_1101001111110000_0101000100000000"; -- -0.1721143126487732
	pesos_i(92) := b"1111111111111111_1111111111111111_1111000111011100_1001100101010000"; -- -0.05522767826914787
	pesos_i(93) := b"1111111111111111_1111111111111111_1110010111001110_0011100100100000"; -- -0.1023220345377922
	pesos_i(94) := b"1111111111111111_1111111111111111_1100111010111101_1010100111000000"; -- -0.19241847097873688
	pesos_i(95) := b"0000000000000000_0000000000000000_0100010010101000_0110111100000000"; -- 0.26819509267807007
	pesos_i(96) := b"1111111111111111_1111111111111111_1111110010010101_1110101101011000"; -- -0.013337412849068642
	pesos_i(97) := b"1111111111111111_1111111111111111_1110001111010111_1100001111000000"; -- -0.10998894274234772
	pesos_i(98) := b"0000000000000000_0000000000000000_0000111010001101_0110100010110000"; -- 0.056845229119062424
	pesos_i(99) := b"0000000000000000_0000000000000000_0000001100001011_1001011111110000"; -- 0.011895652860403061
	pesos_i(100) := b"0000000000000000_0000000000000000_0011001101000110_1010111001000000"; -- 0.2002972513437271
	pesos_i(101) := b"0000000000000000_0000000000000000_0001001101011101_1010001100000000"; -- 0.07564753293991089
	pesos_i(102) := b"0000000000000000_0000000000000000_0000000010010100_0010010111011001"; -- 0.0022605566773563623
	pesos_i(103) := b"1111111111111111_1111111111111111_1111010001011110_0110111010010000"; -- -0.04543408378958702
	pesos_i(104) := b"1111111111111111_1111111111111111_1101000010111010_0011001010000000"; -- -0.18465885519981384
	pesos_i(105) := b"1111111111111111_1111111111111111_1111001010100101_1111001011110000"; -- -0.05215531960129738
	pesos_i(106) := b"1111111111111111_1111111111111111_1110011111010010_1100001110000000"; -- -0.09444025158882141
	pesos_i(107) := b"0000000000000000_0000000000000000_0000011010010010_0110101001011000"; -- 0.025671621784567833
	pesos_i(108) := b"0000000000000000_0000000000000000_0000100110111011_0000010011100000"; -- 0.03800993412733078
	pesos_i(109) := b"1111111111111111_1111111111111111_1100110100000110_0000110000000000"; -- -0.1991264820098877
	pesos_i(110) := b"0000000000000000_0000000000000000_0001101011111100_0101111011100000"; -- 0.10541336983442307
	pesos_i(111) := b"0000000000000000_0000000000000000_0011000110000000_0011010111000000"; -- 0.19336257874965668
	pesos_i(112) := b"0000000000000000_0000000000000000_0011000100101000_1100101111000000"; -- 0.19202874600887299
	pesos_i(113) := b"1111111111111111_1111111111111111_1111101010110001_0000111111101000"; -- -0.02073574624955654
	pesos_i(114) := b"1111111111111111_1111111111111111_1110001000111001_0001010111000000"; -- -0.11631645262241364
	pesos_i(115) := b"1111111111111111_1111111111111111_1011110010010101_1000011010000000"; -- -0.2633434236049652
	pesos_i(116) := b"0000000000000000_0000000000000000_0000001011010011_0001001011000100"; -- 0.011033223010599613
	pesos_i(117) := b"1111111111111111_1111111111111111_1110111010011110_1100111101000000"; -- -0.0678892582654953
	pesos_i(118) := b"1111111111111111_1111111111111111_1101100110100100_1010110011000000"; -- -0.14983101189136505
	pesos_i(119) := b"0000000000000000_0000000000000000_0000101111001000_0000110110000000"; -- 0.04602131247520447
	pesos_i(120) := b"1111111111111111_1111111111111111_1110101001101001_1011010110100000"; -- -0.08432450145483017
	pesos_i(121) := b"0000000000000000_0000000000000000_0011010101111000_0010000101000000"; -- 0.20886428654193878
	pesos_i(122) := b"0000000000000000_0000000000000000_0000010110111001_1101111000100000"; -- 0.022367365658283234
	pesos_i(123) := b"1111111111111111_1111111111111111_1111100111111001_0110110001011000"; -- -0.023537853732705116
	pesos_i(124) := b"1111111111111111_1111111111111111_1111101001110110_0000100100111000"; -- -0.021636413410305977
	pesos_i(125) := b"1111111111111111_1111111111111111_1110001010010010_0001100100000000"; -- -0.11495822668075562
	pesos_i(126) := b"1111111111111111_1111111111111111_1111001101111001_0110111100010000"; -- -0.04892831668257713
	pesos_i(127) := b"0000000000000000_0000000000000000_0011001011001011_1000101000000000"; -- 0.1984182596206665
	pesos_i(128) := b"1111111111111111_1111111111111111_1111111110000101_1101000011110001"; -- -0.0018643771763890982
	pesos_i(129) := b"1111111111111111_1111111111111111_1100101101100000_0101000111000000"; -- -0.2055615335702896
	pesos_i(130) := b"1111111111111111_1111111111111111_1111011001010100_0000011001110000"; -- -0.03778037801384926
	pesos_i(131) := b"1111111111111111_1111111111111111_1111011011110101_0111111100000000"; -- -0.035316526889801025
	pesos_i(132) := b"1111111111111111_1111111111111111_1110100100001100_0011001110100000"; -- -0.08965756744146347
	pesos_i(133) := b"1111111111111111_1111111111111111_1110100000110001_1100000000100000"; -- -0.09299086779356003
	pesos_i(134) := b"0000000000000000_0000000000000000_0100000100000101_1010100000000000"; -- 0.25399255752563477
	pesos_i(135) := b"0000000000000000_0000000000000000_0010100100100111_1111100001000000"; -- 0.160766139626503
	pesos_i(136) := b"1111111111111111_1111111111111111_1100100101111010_1100011110000000"; -- -0.2129702866077423
	pesos_i(137) := b"1111111111111111_1111111111111111_1101110110011100_0001100011000000"; -- -0.1343369036912918
	pesos_i(138) := b"1111111111111111_1111111111111111_1110111100011011_1100110000000000"; -- -0.06598210334777832
	pesos_i(139) := b"0000000000000000_0000000000000000_0011011111111110_0010110011000000"; -- 0.2187221497297287
	pesos_i(140) := b"1111111111111111_1111111111111111_1111101001101010_0010101011111000"; -- -0.021817507222294807
	pesos_i(141) := b"1111111111111111_1111111111111111_1111000101011000_1001100101110000"; -- -0.057241830974817276
	pesos_i(142) := b"0000000000000000_0000000000000000_0000010111101111_1101010100000000"; -- 0.023190796375274658
	pesos_i(143) := b"1111111111111111_1111111111111111_1110000010100011_0000011011100000"; -- -0.12251240760087967
	pesos_i(144) := b"0000000000000000_0000000000000000_0010000111111110_1010000101000000"; -- 0.13279159367084503
	pesos_i(145) := b"0000000000000000_0000000000000000_0010101110101110_0110101000000000"; -- 0.1706300973892212
	pesos_i(146) := b"0000000000000000_0000000000000000_0000011100001110_1011111111100000"; -- 0.027568809688091278
	pesos_i(147) := b"1111111111111111_1111111111111111_1110110010000010_0110011111000000"; -- -0.07613517343997955
	pesos_i(148) := b"0000000000000000_0000000000000000_0001001110101101_0100001011100000"; -- 0.07686250656843185
	pesos_i(149) := b"1111111111111111_1111111111111111_1101111011110100_1101100111000000"; -- -0.12907637655735016
	pesos_i(150) := b"1111111111111111_1111111111111111_1101100000101011_1010001011000000"; -- -0.1555841714143753
	pesos_i(151) := b"1111111111111111_1111111111111111_1111001110000110_0111110110010000"; -- -0.04872908815741539
	pesos_i(152) := b"1111111111111111_1111111111111111_1101110111101010_1010101001000000"; -- -0.133138045668602
	pesos_i(153) := b"1111111111111111_1111111111111111_1011100110110111_1000101100000000"; -- -0.2745431065559387
	pesos_i(154) := b"1111111111111111_1111111111111111_1110101011011000_0101000101100000"; -- -0.0826367512345314
	pesos_i(155) := b"1111111111111111_1111111111111111_1111011110101111_0111110101110000"; -- -0.03247848525643349
	pesos_i(156) := b"0000000000000000_0000000000000000_0110100110101100_0010001100000000"; -- 0.41278284788131714
	pesos_i(157) := b"0000000000000000_0000000000000000_0011110100010011_0100001101000000"; -- 0.23857517540454865
	pesos_i(158) := b"1111111111111111_1111111111111111_1101111001001100_1011010101000000"; -- -0.13164202868938446
	pesos_i(159) := b"0000000000000000_0000000000000000_0001001010101001_1100110001100000"; -- 0.07290341705083847
	pesos_i(160) := b"0000000000000000_0000000000000000_0100111010100100_0101010000000000"; -- 0.30719494819641113
	pesos_i(161) := b"1111111111111111_1111111111111111_1100000100110100_1010000010000000"; -- -0.24529072642326355
	pesos_i(162) := b"0000000000000000_0000000000000000_0110000111000001_0100010010000000"; -- 0.3818552792072296
	pesos_i(163) := b"0000000000000000_0000000000000000_0001100001010010_0001001001000000"; -- 0.09500230848789215
	pesos_i(164) := b"1111111111111111_1111111111111111_1110011011111110_0110111000000000"; -- -0.09768021106719971
	pesos_i(165) := b"0000000000000000_0000000000000000_0001111000100000_0001111000000000"; -- 0.11767756938934326
	pesos_i(166) := b"1111111111111111_1111111111111111_1111000001001101_0111000001010000"; -- -0.061318378895521164
	pesos_i(167) := b"0000000000000000_0000000000000000_0001100010010101_1001111011000000"; -- 0.0960330218076706
	pesos_i(168) := b"1111111111111111_1111111111111111_1110100001101101_0100010111000000"; -- -0.09208263456821442
	pesos_i(169) := b"0000000000000000_0000000000000000_0010001111100011_1000111000000000"; -- 0.1401909589767456
	pesos_i(170) := b"0000000000000000_0000000000000000_0101110101100000_0001000000000000"; -- 0.3647470474243164
	pesos_i(171) := b"0000000000000000_0000000000000000_0010111111010100_1110001001000000"; -- 0.18684209883213043
	pesos_i(172) := b"1111111111111111_1111111111111111_1011000110101111_1100000010000000"; -- -0.30591198801994324
	pesos_i(173) := b"0000000000000000_0000000000000000_0100111000100101_0000100000000000"; -- 0.3052525520324707
	pesos_i(174) := b"1111111111111111_1111111111111111_1100101011110000_0100011000000000"; -- -0.20727121829986572
	pesos_i(175) := b"1111111111111111_1111111111111111_1011100011110011_0001000100000000"; -- -0.2775411009788513
	pesos_i(176) := b"1111111111111111_1111111111111111_1111001101110111_1101001110010000"; -- -0.048952843993902206
	pesos_i(177) := b"0000000000000000_0000000000000000_0010110000100010_1110011100000000"; -- 0.17240756750106812
	pesos_i(178) := b"0000000000000000_0000000000000000_0001101101101101_0011000111000000"; -- 0.10713492333889008
	pesos_i(179) := b"0000000000000000_0000000000000000_0000110100110011_1101110010000000"; -- 0.051572591066360474
	pesos_i(180) := b"1111111111111111_1111111111111111_1111000010011101_0100110000000000"; -- -0.06009984016418457
	pesos_i(181) := b"1111111111111111_1111111111111111_1011010101000100_1101110010000000"; -- -0.291918009519577
	pesos_i(182) := b"1111111111111111_1111111111111111_1110011011111001_1000010000000000"; -- -0.09775519371032715
	pesos_i(183) := b"1111111111111111_1111111111111111_1100001101011100_1000001001000000"; -- -0.236869677901268
	pesos_i(184) := b"1111111111111111_1111111111111111_1110001001110000_1000011100000000"; -- -0.11547046899795532
	pesos_i(185) := b"0000000000000000_0000000000000000_0001001101000011_1110101000000000"; -- 0.07525503635406494
	pesos_i(186) := b"0000000000000000_0000000000000000_0000111110110010_1110010110000000"; -- 0.06132349371910095
	pesos_i(187) := b"0000000000000000_0000000000000000_0110110011111110_0010011110000000"; -- 0.42575308680534363
	pesos_i(188) := b"1111111111111111_1111111111111111_1111111001111101_1010110101110100"; -- -0.005894812755286694
	pesos_i(189) := b"1111111111111111_1111111111111111_1111110111101111_0100001100010100"; -- -0.008067901246249676
	pesos_i(190) := b"0000000000000000_0000000000000000_0010010100110110_0101010011000000"; -- 0.14536027610301971
	pesos_i(191) := b"0000000000000000_0000000000000000_0000001010101010_1101011110111100"; -- 0.010419352911412716
	pesos_i(192) := b"1111111111111111_1111111111111111_1101100100101011_0100111000000000"; -- -0.15168297290802002
	pesos_i(193) := b"1111111111111111_1111111111111111_1111011010010110_0111000110000000"; -- -0.03676691651344299
	pesos_i(194) := b"0000000000000000_0000000000000000_0001100111001111_0000101100100000"; -- 0.10081548243761063
	pesos_i(195) := b"0000000000000000_0000000000000000_0000000011001000_1111001000101010"; -- 0.003066191915422678
	pesos_i(196) := b"1111111111111111_1111111111111111_1010110110011101_1000111100000000"; -- -0.3218145966529846
	pesos_i(197) := b"0000000000000000_0000000000000000_0001111010001100_0111011000100000"; -- 0.11933077126741409
	pesos_i(198) := b"0000000000000000_0000000000000000_0011100001101111_0001010001000000"; -- 0.2204449325799942
	pesos_i(199) := b"1111111111111111_1111111111111111_1010001000101111_0111100100000000"; -- -0.3664631247520447
	pesos_i(200) := b"1111111111111111_1111111111111111_1101010010101011_0001010010000000"; -- -0.1692645251750946
	pesos_i(201) := b"0000000000000000_0000000000000000_0000111001100101_1111110101110000"; -- 0.05624374374747276
	pesos_i(202) := b"0000000000000000_0000000000000000_0011011101110000_1010010011000000"; -- 0.21656255424022675
	pesos_i(203) := b"0000000000000000_0000000000000000_0100001000110011_1101110010000000"; -- 0.2586038410663605
	pesos_i(204) := b"1111111111111111_1111111111111111_1110001000101010_1110111110100000"; -- -0.1165323480963707
	pesos_i(205) := b"1111111111111111_1111111111111111_1101100110001101_1100011111000000"; -- -0.15018035471439362
	pesos_i(206) := b"1111111111111111_1111111111111111_1101011011011111_1110001111000000"; -- -0.1606462150812149
	pesos_i(207) := b"1111111111111111_1111111111111111_1110011111010000_0101100011100000"; -- -0.09447712451219559
	pesos_i(208) := b"1111111111111111_1111111111111111_1101001010100001_1011010000000000"; -- -0.17722010612487793
	pesos_i(209) := b"0000000000000000_0000000000000000_0101111100101000_1110110100000000"; -- 0.37171822786331177
	pesos_i(210) := b"0000000000000000_0000000000000000_0011000111010010_0001010000000000"; -- 0.1946117877960205
	pesos_i(211) := b"1111111111111111_1111111111111111_1110111100101111_0000110010000000"; -- -0.06568834185600281
	pesos_i(212) := b"1111111111111111_1111111111111111_1010101110001110_1100001110000000"; -- -0.3298528492450714
	pesos_i(213) := b"1111111111111111_1111111111111111_1110001000011110_1000010000100000"; -- -0.11672186106443405
	pesos_i(214) := b"1111111111111111_1111111111111111_1011001100011001_0011110000000000"; -- -0.300396203994751
	pesos_i(215) := b"1111111111111111_1111111111111111_1111010011001110_1000101101110000"; -- -0.04372337833046913
	pesos_i(216) := b"0000000000000000_0000000000000000_0000001111000111_0011100100100000"; -- 0.014758653938770294
	pesos_i(217) := b"0000000000000000_0000000000000000_0010110110010000_1010011000000000"; -- 0.17798840999603271
	pesos_i(218) := b"1111111111111111_1111111111111111_1001001000110010_0010101010000000"; -- -0.42892202734947205
	pesos_i(219) := b"1111111111111111_1111111111111111_1011000010000001_1101000100000000"; -- -0.31051915884017944
	pesos_i(220) := b"1111111111111111_1111111111111111_1110000111000000_1001110010000000"; -- -0.11815473437309265
	pesos_i(221) := b"1111111111111111_1111111111111111_1110100000000100_0001010011000000"; -- -0.09368772804737091
	pesos_i(222) := b"0000000000000000_0000000000000000_0011011101001011_1001111100000000"; -- 0.2159976363182068
	pesos_i(223) := b"1111111111111111_1111111111111111_1111010011111010_1110111111100000"; -- -0.0430460050702095
	pesos_i(224) := b"0000000000000000_0000000000000000_0001010011100001_0010010010100000"; -- 0.0815604105591774
	pesos_i(225) := b"0000000000000000_0000000000000000_0001100010000111_0110101011000000"; -- 0.09581629931926727
	pesos_i(226) := b"0000000000000000_0000000000000000_0000011011011110_1011010001011000"; -- 0.026835700497031212
	pesos_i(227) := b"0000000000000000_0000000000000000_0001001100000001_1010111000000000"; -- 0.07424437999725342
	pesos_i(228) := b"1111111111111111_1111111111111111_1110100000001110_0011011101000000"; -- -0.09353308379650116
	pesos_i(229) := b"0000000000000000_0000000000000000_0010110100001000_1000110011000000"; -- 0.17591170966625214
	pesos_i(230) := b"1111111111111111_1111111111111111_1111001100011001_1011010011000000"; -- -0.05038900673389435
	pesos_i(231) := b"0000000000000000_0000000000000000_0000100011000000_0110000110010000"; -- 0.0341855026781559
	pesos_i(232) := b"1111111111111111_1111111111111111_1111011011001001_0111000000100000"; -- -0.03598880022764206
	pesos_i(233) := b"0000000000000000_0000000000000000_0011100111001110_0001110100000000"; -- 0.2258012890815735
	pesos_i(234) := b"1111111111111111_1111111111111111_1110011110011001_0010010010100000"; -- -0.0953194722533226
	pesos_i(235) := b"0000000000000000_0000000000000000_0010001000010111_1100011010000000"; -- 0.13317528367042542
	pesos_i(236) := b"0000000000000000_0000000000000000_0010011001011000_1000101010000000"; -- 0.1497885286808014
	pesos_i(237) := b"1111111111111111_1111111111111111_1100110111101011_0110010111000000"; -- -0.1956268697977066
	pesos_i(238) := b"1111111111111111_1111111111111111_1111101010110111_1101111101011000"; -- -0.020631829276680946
	pesos_i(239) := b"0000000000000000_0000000000000000_0000011010110110_0111101100000000"; -- 0.026221930980682373
	pesos_i(240) := b"1111111111111111_1111111111111111_1010010101110100_0000001100000000"; -- -0.3536985516548157
	pesos_i(241) := b"1111111111111111_1111111111111111_1011100101011101_0001100010000000"; -- -0.2759232223033905
	pesos_i(242) := b"0000000000000000_0000000000000000_0100001111111011_1110011110000000"; -- 0.265562504529953
	pesos_i(243) := b"1111111111111111_1111111111111111_1001001000101011_0111100000000000"; -- -0.42902421951293945
	pesos_i(244) := b"1111111111111111_1111111111111111_1010011100101001_0100010010000000"; -- -0.3470265567302704
	pesos_i(245) := b"0000000000000000_0000000000000000_0011110101110101_1100000010000000"; -- 0.24007800221443176
	pesos_i(246) := b"1111111111111111_1111111111111111_1101111111001111_0011010011000000"; -- -0.1257445365190506
	pesos_i(247) := b"1111111111111111_1111111111111111_1101100100010100_1001000110000000"; -- -0.15202990174293518
	pesos_i(248) := b"0000000000000000_0000000000000000_0001101001110000_0011111101100000"; -- 0.10327526181936264
	pesos_i(249) := b"0000000000000000_0000000000000000_0011000101110011_0011011110000000"; -- 0.19316431879997253
	pesos_i(250) := b"1111111111111111_1111111111111111_1111101101001110_1100100000111000"; -- -0.018329130485653877
	pesos_i(251) := b"0000000000000000_0000000000000000_0010000001001110_1000101010000000"; -- 0.1261984407901764
	pesos_i(252) := b"0000000000000000_0000000000000000_0100001100011011_1100100010000000"; -- 0.26214268803596497
	pesos_i(253) := b"1111111111111111_1111111111111111_1110000100111101_0110001100000000"; -- -0.12015706300735474
	pesos_i(254) := b"1111111111111111_1111111111111111_1101010100001000_1101001010000000"; -- -0.16783413290977478
	pesos_i(255) := b"0000000000000000_0000000000000000_0000000110010000_1001101110100110"; -- 0.006112792994827032
	pesos_i(256) := b"0000000000000000_0000000000000000_0101110110101001_1001011100000000"; -- 0.3658689856529236
	pesos_i(257) := b"1111111111111111_1111111111111111_1000010100100110_1001100010000000"; -- -0.47987982630729675
	pesos_i(258) := b"0000000000000000_0000000000000000_0010011100000101_0100101011000000"; -- 0.15242449939250946
	pesos_i(259) := b"0000000000000000_0000000000000000_0001011001101011_0010011101100000"; -- 0.08757253736257553
	pesos_i(260) := b"1111111111111111_1111111111111111_1010011110010011_0101000010000000"; -- -0.3454084098339081
	pesos_i(261) := b"0000000000000000_0000000000000000_0000010111010011_1111100110001000"; -- 0.02276572771370411
	pesos_i(262) := b"0000000000000000_0000000000000000_1001100000101011_1001010100000000"; -- 0.594415009021759
	pesos_i(263) := b"1111111111111111_1111111111111111_1111111000000100_0110011101110010"; -- -0.007745299022644758
	pesos_i(264) := b"1111111111111111_1111111111111111_0100101010100110_1001101100000000"; -- -0.7083953022956848
	pesos_i(265) := b"1111111111111111_1111111111111111_1110111111001001_0101000010000000"; -- -0.06333443522453308
	pesos_i(266) := b"1111111111111111_1111111111111111_1100000010110110_0001000011000000"; -- -0.247221902012825
	pesos_i(267) := b"0000000000000000_0000000000000000_0111011011001110_1001010000000000"; -- 0.46408963203430176
	pesos_i(268) := b"0000000000000000_0000000000000000_0010011011001011_0101001111000000"; -- 0.15154002606868744
	pesos_i(269) := b"0000000000000000_0000000000000000_0101110011110010_1110110100000000"; -- 0.36308175325393677
	pesos_i(270) := b"0000000000000000_0000000000000000_1011110101011000_1101000000000000"; -- 0.7396364212036133
	pesos_i(271) := b"1111111111111111_1111111111111111_1001000110111000_1011010110000000"; -- -0.43077531456947327
	pesos_i(272) := b"0000000000000000_0000000000000000_0011000111001010_1010110000000000"; -- 0.19449877738952637
	pesos_i(273) := b"0000000000000000_0000000000000000_1111101011101010_1001100100000000"; -- 0.9801421761512756
	pesos_i(274) := b"0000000000000000_0000000000000000_0000111111110011_1100010101100000"; -- 0.06231340020895004
	pesos_i(275) := b"0000000000000000_0000000000000000_0110111000000110_0010001010000000"; -- 0.42978110909461975
	pesos_i(276) := b"0000000000000000_0000000000000000_1001111111100000_0010100000000000"; -- 0.624514102935791
	pesos_i(277) := b"1111111111111111_1111111111111111_1111011001111100_0111101101000000"; -- -0.03716306388378143
	pesos_i(278) := b"1111111111111111_1111111111111111_1111101000111010_0110010100110000"; -- -0.02254645898938179
	pesos_i(279) := b"1111111111111111_1111111111111111_1010111001011100_0011011100000000"; -- -0.31890541315078735
	pesos_i(280) := b"1111111111111111_1111111111111111_0011011100111100_0000010000000000"; -- -0.7842404842376709
	pesos_i(281) := b"1111111111111111_1111111111111111_1010100111001000_0101010000000000"; -- -0.33678698539733887
	pesos_i(282) := b"1111111111111111_1111111111111111_1111101111010010_0011001100010000"; -- -0.016323860734701157
	pesos_i(283) := b"0000000000000000_0000000000000000_0001110001110101_1001111110000000"; -- 0.11116978526115417
	pesos_i(284) := b"0000000000000000_0000000000000000_1001001110100001_0100001000000000"; -- 0.5766793489456177
	pesos_i(285) := b"0000000000000000_0000000000000000_0100011011100110_0011001000000000"; -- 0.27695000171661377
	pesos_i(286) := b"1111111111111111_1111111111111111_0101001110001101_1111100100000000"; -- -0.6736149191856384
	pesos_i(287) := b"0000000000000000_0000000000000000_0011110100001111_1101000110000000"; -- 0.23852261900901794
	pesos_i(288) := b"0000000000000000_0000000000000000_0010011001000100_0101110110000000"; -- 0.1494806706905365
	pesos_i(289) := b"1111111111111111_1111111111111111_1111000010101110_0101101111010000"; -- -0.05983949825167656
	pesos_i(290) := b"0000000000000000_0000000000000000_1000000001001000_0001100100000000"; -- 0.5011001229286194
	pesos_i(291) := b"0000000000000000_0000000000000000_0101100011111110_1101100010000000"; -- 0.34763863682746887
	pesos_i(292) := b"1111111111111111_1111111111111111_1100101000000101_0001111000000000"; -- -0.21085941791534424
	pesos_i(293) := b"0000000000000000_0000000000000000_1000010101101010_0101100100000000"; -- 0.52115398645401
	pesos_i(294) := b"1111111111111111_1111111111111111_1101000011001011_0000011001000000"; -- -0.18440209329128265
	pesos_i(295) := b"1111111111111111_1111111111111111_1010111010010101_0111100100000000"; -- -0.3180317282676697
	pesos_i(296) := b"0000000000000000_0000000000000000_0001100101000001_0101111101000000"; -- 0.09865374863147736
	pesos_i(297) := b"0000000000000000_0000000000000000_1010000011110111_0001110100000000"; -- 0.628770649433136
	pesos_i(298) := b"0000000000000000_0000000000000000_0011100100000011_1010110011000000"; -- 0.22271232306957245
	pesos_i(299) := b"0000000000000000_0000000000000000_0000011000001111_0100101011101000"; -- 0.023670846596360207
	pesos_i(300) := b"1111111111111111_1111111111111111_1011000101011111_0110000000000000"; -- -0.30713844299316406
	pesos_i(301) := b"0000000000000000_0000000000000000_0111110000010101_1110100010000000"; -- 0.4847092926502228
	pesos_i(302) := b"1111111111111111_1111111111111111_0111010111010000_0000111100000000"; -- -0.5397940278053284
	pesos_i(303) := b"1111111111111111_1111111111111111_1101101011110010_1101001101000000"; -- -0.1447322815656662
	pesos_i(304) := b"1111111111111111_1111111111111111_1100011111101001_1001110111000000"; -- -0.21909154951572418
	pesos_i(305) := b"0000000000000000_0000000000000000_0100011001101110_0011110110000000"; -- 0.2751196324825287
	pesos_i(306) := b"1111111111111111_1111111111111111_1011001101011111_1011101100000000"; -- -0.2993205189704895
	pesos_i(307) := b"0000000000000000_0000000000000000_0111100011010110_1001101110000000"; -- 0.4720246493816376
	pesos_i(308) := b"1111111111111111_1111111111111111_0111101100111110_1011110000000000"; -- -0.5185739994049072
	pesos_i(309) := b"1111111111111111_1111111111111111_0111111101001010_0111100100000000"; -- -0.5027698874473572
	pesos_i(310) := b"0000000000000000_0000000000000000_0110101101011101_0001011100000000"; -- 0.41938918828964233
	pesos_i(311) := b"1111111111111111_1111111111111111_1101111111010110_1110000001000000"; -- -0.12562750279903412
	pesos_i(312) := b"1111111111111111_1111111111111111_1011110011101001_0100100110000000"; -- -0.2620653212070465
	pesos_i(313) := b"0000000000000000_0000000000000000_0000001101000101_0000101011101100"; -- 0.012772257439792156
	pesos_i(314) := b"1111111111111111_1111111111111111_1101110110011111_1000000111000000"; -- -0.1342848688364029
	pesos_i(315) := b"0000000000000000_0000000000000000_1000010010101001_0010000100000000"; -- 0.5182057023048401
	pesos_i(316) := b"1111111111111111_1111111111111111_1101010011110111_1110011011000000"; -- -0.16809232532978058
	pesos_i(317) := b"0000000000000000_0000000000000000_0011011011101011_0000000101000000"; -- 0.21452338993549347
	pesos_i(318) := b"0000000000000000_0000000000000000_0100010110110100_1111010110000000"; -- 0.27229246497154236
	pesos_i(319) := b"0000000000000000_0000000000000000_1010000000011010_1101111100000000"; -- 0.6254100203514099
	pesos_i(320) := b"1111111111111111_1111111111111111_1111011101010010_0111001100100000"; -- -0.03389816731214523
	pesos_i(321) := b"1111111111111111_1111111111111111_1101100100111111_0111001100000000"; -- -0.15137559175491333
	pesos_i(322) := b"0000000000000000_0000000000000000_0110001000000001_1011000010000000"; -- 0.38283827900886536
	pesos_i(323) := b"0000000000000000_0000000000000000_0011000010000111_1110010001000000"; -- 0.18957354128360748
	pesos_i(324) := b"1111111111111111_1111111111111111_1000100110111110_0100000100000000"; -- -0.4619407057762146
	pesos_i(325) := b"0000000000000000_0000000000000000_1000100011000001_1100000000000000"; -- 0.5342063903808594
	pesos_i(326) := b"0000000000000000_0000000000000000_0010001110111001_0001100101000000"; -- 0.13954313099384308
	pesos_i(327) := b"1111111111111111_1111111111111111_0110000001000011_0101101000000000"; -- -0.6239722967147827
	pesos_i(328) := b"0000000000000000_0000000000000000_0100111100011111_0101000010000000"; -- 0.3090715706348419
	pesos_i(329) := b"1111111111111111_1111111111111111_1011111000010110_1100100100000000"; -- -0.25746482610702515
	pesos_i(330) := b"0000000000000000_0000000000000000_0001110000000011_1000011101000000"; -- 0.10942883789539337
	pesos_i(331) := b"1111111111111111_1111111111111111_1110111010111101_0111111001000000"; -- -0.0674210637807846
	pesos_i(332) := b"1111111111111111_1111111111111111_1100001010000011_0111101000000000"; -- -0.2401813268661499
	pesos_i(333) := b"0000000000000000_0000000000000000_0001101100111010_1011111010000000"; -- 0.10636511445045471
	pesos_i(334) := b"1111111111111111_1111111111111111_1100010111101001_1110111000000000"; -- -0.22689926624298096
	pesos_i(335) := b"1111111111111111_1111111111111111_1111101011100011_1001110101001000"; -- -0.01996438018977642
	pesos_i(336) := b"0000000000000000_0000000000000000_0010011110100111_0100001011000000"; -- 0.15489594638347626
	pesos_i(337) := b"0000000000000000_0000000000000000_0011010110000011_1010000000000000"; -- 0.20903968811035156
	pesos_i(338) := b"0000000000000000_0000000000000000_0101011111101101_0110101010000000"; -- 0.3434664309024811
	pesos_i(339) := b"0000000000000000_0000000000000000_1001010111111100_1110011000000000"; -- 0.5858901739120483
	pesos_i(340) := b"1111111111111111_1111111111111111_0001100100100000_0110110100000000"; -- -0.9018489718437195
	pesos_i(341) := b"1111111111111111_1111111111111111_0010111011100101_1111100000000000"; -- -0.8168034553527832
	pesos_i(342) := b"1111111111111111_1111111111111111_0101101110000100_0001011100000000"; -- -0.6425157189369202
	pesos_i(343) := b"1111111111111111_1111111111111111_0110001111111010_1100011100000000"; -- -0.6094546914100647
	pesos_i(344) := b"1111111111111111_1111111111111111_1110001001000111_1111001101100000"; -- -0.11608961969614029
	pesos_i(345) := b"0000000000000000_0000000000000000_0000110110110011_1111001000110000"; -- 0.05352700874209404
	pesos_i(346) := b"1111111111111111_1111111111111111_0110110100011100_1111101100000000"; -- -0.5737765431404114
	pesos_i(347) := b"1111111111111111_1111111111111111_1011101010010101_1000000100000000"; -- -0.2711562514305115
	pesos_i(348) := b"0000000000000000_0000000000000000_0100010011111011_1001100100000000"; -- 0.26946407556533813
	pesos_i(349) := b"1111111111111111_1111111111111111_1000001100100100_0110111100000000"; -- -0.48772531747817993
	pesos_i(350) := b"0000000000000000_0000000000000000_0011100111000110_1001101110000000"; -- 0.22568675875663757
	pesos_i(351) := b"0000000000000000_0000000000000000_0001011101110001_0010010011100000"; -- 0.09157019108533859
	pesos_i(352) := b"0000000000000000_0000000000000000_0000111100011011_1101111001010000"; -- 0.05901898816227913
	pesos_i(353) := b"0000000000000000_0000000000000000_0000000101011100_1000000100000000"; -- 0.005317747592926025
	pesos_i(354) := b"1111111111111111_1111111111111111_1010111110100100_1101001100000000"; -- -0.3138912320137024
	pesos_i(355) := b"1111111111111111_1111111111111111_1100101011010011_0000001010000000"; -- -0.20771774649620056
	pesos_i(356) := b"1111111111111111_1111111111111111_1100010111110010_1001111100000000"; -- -0.2267666459083557
	pesos_i(357) := b"0000000000000000_0000000000000000_0010001111110110_0000000011000000"; -- 0.14047245681285858
	pesos_i(358) := b"1111111111111111_1111111111111111_1010001110100011_1100111010000000"; -- -0.3607817590236664
	pesos_i(359) := b"0000000000000000_0000000000000000_0000100011101100_1011000100100000"; -- 0.03486163169145584
	pesos_i(360) := b"1111111111111111_1111111111111111_1100011110010001_0010101100000000"; -- -0.22044116258621216
	pesos_i(361) := b"1111111111111111_1111111111111111_1011001110110000_1100000010000000"; -- -0.29808422923088074
	pesos_i(362) := b"0000000000000000_0000000000000000_0000101100011111_0111100010110000"; -- 0.04344896599650383
	pesos_i(363) := b"0000000000000000_0000000000000000_0101110000000010_1111011000000000"; -- 0.35942018032073975
	pesos_i(364) := b"0000000000000000_0000000000000000_0011111110100100_0011101100000000"; -- 0.24859970808029175
	pesos_i(365) := b"1111111111111111_1111111111111111_1110001010111110_0011000001100000"; -- -0.11428544670343399
	pesos_i(366) := b"0000000000000000_0000000000000000_0111011010001110_1001110110000000"; -- 0.4631136357784271
	pesos_i(367) := b"0000000000000000_0000000000000000_0000010110100000_1010000000110000"; -- 0.021982204169034958
	pesos_i(368) := b"1111111111111111_1111111111111111_1001011111110101_0101011010000000"; -- -0.40641269087791443
	pesos_i(369) := b"1111111111111111_1111111111111111_1110111000100001_0001111110100000"; -- -0.06980707496404648
	pesos_i(370) := b"0000000000000000_0000000000000000_1000000110010111_1100011000000000"; -- 0.506222128868103
	pesos_i(371) := b"1111111111111111_1111111111111111_0100111100000111_0011111100000000"; -- -0.6912956833839417
	pesos_i(372) := b"1111111111111111_1111111111111111_0010001111100101_1010101000000000"; -- -0.8597768545150757
	pesos_i(373) := b"0000000000000000_0000000000000000_0111010010001111_1111001010000000"; -- 0.45532146096229553
	pesos_i(374) := b"0000000000000000_0000000000000000_0010000101000010_0001101101000000"; -- 0.12991495430469513
	pesos_i(375) := b"1111111111111111_1111111111111111_1111101111011010_0011000000110000"; -- -0.016201961785554886
	pesos_i(376) := b"0000000000000000_0000000000000000_0110101100111110_1000111010000000"; -- 0.4189232885837555
	pesos_i(377) := b"0000000000000000_0000000000000000_1100100111011010_0010001100000000"; -- 0.7884847521781921
	pesos_i(378) := b"0000000000000000_0000000000000000_0001101010000101_1010110011100000"; -- 0.10360222309827805
	pesos_i(379) := b"1111111111111111_1111111111111111_1000011000101110_0101001100000000"; -- -0.47585564851760864
	pesos_i(380) := b"0000000000000000_0000000000000000_0011111000010011_1101100001000000"; -- 0.24249030649662018
	pesos_i(381) := b"1111111111111111_1111111111111111_1110000110100100_1001110101000000"; -- -0.11858193576335907
	pesos_i(382) := b"1111111111111111_1111111111111111_1111100010111010_0001110100010000"; -- -0.028410132974386215
	pesos_i(383) := b"0000000000000000_0000000000000000_0101110111110111_0010100000000000"; -- 0.3670525550842285
	pesos_i(384) := b"0000000000000000_0000000000000000_1100011100000100_0110000000000000"; -- 0.7774105072021484
	pesos_i(385) := b"1111111111111111_1111111111111110_1110111111001011_1001011000000000"; -- -1.0632997751235962
	pesos_i(386) := b"0000000000000000_0000000000000000_0100100101101001_0011001010000000"; -- 0.28676143288612366
	pesos_i(387) := b"1111111111111111_1111111111111111_1110011111110011_0111010001000000"; -- -0.09394143521785736
	pesos_i(388) := b"1111111111111111_1111111111111111_0101010000101010_0110111000000000"; -- -0.6712275743484497
	pesos_i(389) := b"0000000000000000_0000000000000000_0111101100101110_0111001000000000"; -- 0.4811774492263794
	pesos_i(390) := b"0000000000000000_0000000000000001_0000100001010101_0010001000000000"; -- 1.0325490236282349
	pesos_i(391) := b"0000000000000000_0000000000000000_0010110000111100_1000001111000000"; -- 0.17279838025569916
	pesos_i(392) := b"1111111111111111_1111111111111110_1111001110000000_0010100000000000"; -- -1.048825740814209
	pesos_i(393) := b"1111111111111111_1111111111111111_0111100011000111_0010000000000000"; -- -0.5282115936279297
	pesos_i(394) := b"1111111111111111_1111111111111111_1000010111000010_1111101110000000"; -- -0.477493554353714
	pesos_i(395) := b"0000000000000000_0000000000000000_1100001111000111_0110111100000000"; -- 0.7647618651390076
	pesos_i(396) := b"0000000000000000_0000000000000000_0000001100110110_0111000101000000"; -- 0.012549474835395813
	pesos_i(397) := b"1111111111111111_1111111111111111_1111110100100101_1101100000100100"; -- -0.011141291819512844
	pesos_i(398) := b"0000000000000000_0000000000000000_1001001001100011_1010110000000000"; -- 0.5718333721160889
	pesos_i(399) := b"1111111111111111_1111111111111111_0111100011100100_0010101000000000"; -- -0.5277684926986694
	pesos_i(400) := b"0000000000000000_0000000000000000_0011001110100110_0001111011000000"; -- 0.20175354182720184
	pesos_i(401) := b"0000000000000000_0000000000000001_0011000100101001_1000100000000000"; -- 1.192039966583252
	pesos_i(402) := b"0000000000000000_0000000000000000_0000101111000001_0001111101110000"; -- 0.045915570110082626
	pesos_i(403) := b"0000000000000000_0000000000000000_1010100000110100_1101110000000000"; -- 0.6570565700531006
	pesos_i(404) := b"0000000000000000_0000000000000000_1001110110010100_0011101100000000"; -- 0.6155430674552917
	pesos_i(405) := b"1111111111111111_1111111111111111_1101000000011101_1100000100000000"; -- -0.18704599142074585
	pesos_i(406) := b"0000000000000000_0000000000000000_0001100110101101_1000101101000000"; -- 0.10030432045459747
	pesos_i(407) := b"1111111111111111_1111111111111111_1000001110111100_1111001110000000"; -- -0.4853980839252472
	pesos_i(408) := b"1111111111111111_1111111111111111_0010010110011000_0110000100000000"; -- -0.8531436324119568
	pesos_i(409) := b"1111111111111111_1111111111111111_0010111101010010_0000101000000000"; -- -0.8151544332504272
	pesos_i(410) := b"0000000000000000_0000000000000000_0011110010100000_1100100000000000"; -- 0.23682832717895508
	pesos_i(411) := b"0000000000000000_0000000000000000_0000110000000001_1101100010010000"; -- 0.04690316691994667
	pesos_i(412) := b"0000000000000000_0000000000000000_1110000000001000_0111110000000000"; -- 0.8751294612884521
	pesos_i(413) := b"0000000000000000_0000000000000000_0100101100000111_1010001100000000"; -- 0.2930852770805359
	pesos_i(414) := b"1111111111111111_1111111111111111_0110101011000011_0110010100000000"; -- -0.5829560160636902
	pesos_i(415) := b"0000000000000000_0000000000000000_0100001101101101_1110000010000000"; -- 0.2633953392505646
	pesos_i(416) := b"0000000000000000_0000000000000000_0111111011111100_0011001100000000"; -- 0.49603575468063354
	pesos_i(417) := b"1111111111111111_1111111111111111_1000011100100011_0110001010000000"; -- -0.4721163213253021
	pesos_i(418) := b"0000000000000000_0000000000000000_1100100010000101_1001001100000000"; -- 0.7832881808280945
	pesos_i(419) := b"0000000000000000_0000000000000000_0110010110110001_0011100110000000"; -- 0.3972354829311371
	pesos_i(420) := b"1111111111111111_1111111111111111_1001111111101110_0001101000000000"; -- -0.37527310848236084
	pesos_i(421) := b"0000000000000000_0000000000000000_1011111101111010_0000010000000000"; -- 0.7479555606842041
	pesos_i(422) := b"1111111111111111_1111111111111111_1110011101010001_1010000010100000"; -- -0.09641071408987045
	pesos_i(423) := b"1111111111111111_1111111111111111_1011100100011110_1001010110000000"; -- -0.2768770754337311
	pesos_i(424) := b"0000000000000000_0000000000000000_0001101010010010_0001101110100000"; -- 0.10379192978143692
	pesos_i(425) := b"0000000000000000_0000000000000001_0001001011010001_1011110000000000"; -- 1.0735127925872803
	pesos_i(426) := b"0000000000000000_0000000000000000_1001101001001011_1100010100000000"; -- 0.6027186512947083
	pesos_i(427) := b"0000000000000000_0000000000000000_0011001010101100_1101000000000000"; -- 0.19794940948486328
	pesos_i(428) := b"1111111111111111_1111111111111111_1000100101010100_0101100110000000"; -- -0.4635566771030426
	pesos_i(429) := b"0000000000000000_0000000000000000_1101000110011001_1111100000000000"; -- 0.8187556266784668
	pesos_i(430) := b"1111111111111111_1111111111111111_0000001011111101_0110010100000000"; -- -0.9883210062980652
	pesos_i(431) := b"1111111111111111_1111111111111111_0111000000100011_0100000100000000"; -- -0.5619620680809021
	pesos_i(432) := b"0000000000000000_0000000000000000_0010011001010100_0110111111000000"; -- 0.14972589910030365
	pesos_i(433) := b"0000000000000000_0000000000000000_0011101001110001_0010011101000000"; -- 0.22828908264636993
	pesos_i(434) := b"1111111111111111_1111111111111111_1001011101010100_0000111010000000"; -- -0.40887364745140076
	pesos_i(435) := b"0000000000000000_0000000000000000_1100010010101100_0001110000000000"; -- 0.7682511806488037
	pesos_i(436) := b"1111111111111111_1111111111111111_0010001001101011_0010110100000000"; -- -0.8655521273612976
	pesos_i(437) := b"1111111111111111_1111111111111111_0010001111101100_1011000000000000"; -- -0.8596696853637695
	pesos_i(438) := b"0000000000000000_0000000000000000_1011001110010100_1110110000000000"; -- 0.701491117477417
	pesos_i(439) := b"1111111111111111_1111111111111111_1001100001000100_1110100000000000"; -- -0.4051985740661621
	pesos_i(440) := b"1111111111111111_1111111111111111_0101001010111100_1111011100000000"; -- -0.6768041253089905
	pesos_i(441) := b"1111111111111111_1111111111111111_1111110010000101_0011001001010000"; -- -0.013592582195997238
	pesos_i(442) := b"1111111111111111_1111111111111111_1001110000110011_1000100110000000"; -- -0.3898386061191559
	pesos_i(443) := b"0000000000000000_0000000000000001_0010000011110101_1100010000000000"; -- 1.1287500858306885
	pesos_i(444) := b"1111111111111111_1111111111111111_1010000000010101_0000010110000000"; -- -0.37467923760414124
	pesos_i(445) := b"1111111111111111_1111111111111111_1111100111010111_1001001011011000"; -- -0.024054357782006264
	pesos_i(446) := b"0000000000000000_0000000000000000_0100000010001010_1010100100000000"; -- 0.25211578607559204
	pesos_i(447) := b"0000000000000000_0000000000000000_1011101100111101_0001011000000000"; -- 0.7314008474349976
	pesos_i(448) := b"1111111111111111_1111111111111111_1110011100110010_1001011000100000"; -- -0.0968843623995781
	pesos_i(449) := b"1111111111111111_1111111111111111_1111110001101001_0110111100000000"; -- -0.014016211032867432
	pesos_i(450) := b"0000000000000000_0000000000000000_0100111101101101_0110100000000000"; -- 0.31026315689086914
	pesos_i(451) := b"0000000000000000_0000000000000000_0011011111001110_0000101111000000"; -- 0.2179877609014511
	pesos_i(452) := b"1111111111111111_1111111111111111_1000100000000111_0011000000000000"; -- -0.4686403274536133
	pesos_i(453) := b"0000000000000000_0000000000000000_1111101100110011_0101110100000000"; -- 0.9812524914741516
	pesos_i(454) := b"1111111111111111_1111111111111111_0111001011010010_1100001100000000"; -- -0.5514715313911438
	pesos_i(455) := b"1111111111111111_1111111111111111_0011100110010011_1100010000000000"; -- -0.7750890254974365
	pesos_i(456) := b"0000000000000000_0000000000000000_0000000111110000_1101110110011010"; -- 0.007581567857414484
	pesos_i(457) := b"1111111111111111_1111111111111111_0111110001000010_0101001100000000"; -- -0.5146129727363586
	pesos_i(458) := b"1111111111111111_1111111111111111_1101101100110001_0111001001000000"; -- -0.1437767595052719
	pesos_i(459) := b"0000000000000000_0000000000000000_0100100111110011_0010010100000000"; -- 0.2888663411140442
	pesos_i(460) := b"1111111111111111_1111111111111111_1000111000110101_1000010010000000"; -- -0.44449588656425476
	pesos_i(461) := b"0000000000000000_0000000000000000_0000100010111110_0000000010010000"; -- 0.034149203449487686
	pesos_i(462) := b"1111111111111111_1111111111111111_0110010101000100_0000111000000000"; -- -0.6044303178787231
	pesos_i(463) := b"1111111111111111_1111111111111111_1001010110001001_0011010110000000"; -- -0.415875107049942
	pesos_i(464) := b"1111111111111111_1111111111111111_1010001001110001_1001011110000000"; -- -0.36545422673225403
	pesos_i(465) := b"0000000000000000_0000000000000000_1100010010101010_1100010000000000"; -- 0.768230676651001
	pesos_i(466) := b"0000000000000000_0000000000000000_0101010010110000_1010110100000000"; -- 0.33082085847854614
	pesos_i(467) := b"0000000000000000_0000000000000000_0000110111000001_1110110000010000"; -- 0.05374026671051979
	pesos_i(468) := b"1111111111111111_1111111111111110_1100000010100101_0100100000000000"; -- -1.2474780082702637
	pesos_i(469) := b"1111111111111111_1111111111111111_0100011011011101_0110111100000000"; -- -0.7231836915016174
	pesos_i(470) := b"1111111111111111_1111111111111110_1111110001111011_0011110000000000"; -- -1.013744592666626
	pesos_i(471) := b"1111111111111111_1111111111111111_0101011010111100_1011010100000000"; -- -0.6611830592155457
	pesos_i(472) := b"1111111111111111_1111111111111111_1101011010110111_0001001110000000"; -- -0.16126897931098938
	pesos_i(473) := b"1111111111111111_1111111111111111_1110100111100010_0001000011000000"; -- -0.08639426529407501
	pesos_i(474) := b"1111111111111111_1111111111111111_0001000011111101_1111011000000000"; -- -0.9336248636245728
	pesos_i(475) := b"1111111111111111_1111111111111111_1110111001001100_1010010010100000"; -- -0.06914301961660385
	pesos_i(476) := b"0000000000000000_0000000000000000_0101000111101110_1100110100000000"; -- 0.32005006074905396
	pesos_i(477) := b"1111111111111111_1111111111111111_0011011100011100_1000001000000000"; -- -0.7847212553024292
	pesos_i(478) := b"0000000000000000_0000000000000000_0100111000001101_1001010100000000"; -- 0.30489474534988403
	pesos_i(479) := b"0000000000000000_0000000000000000_1010010110110111_0100101000000000"; -- 0.6473280191421509
	pesos_i(480) := b"0000000000000000_0000000000000000_0000001011111011_0110010001010000"; -- 0.011648435145616531
	pesos_i(481) := b"1111111111111111_1111111111111111_1101101011111010_0001101101000000"; -- -0.14462117850780487
	pesos_i(482) := b"0000000000000000_0000000000000000_0000000100110001_0110100011011100"; -- 0.0046601807698607445
	pesos_i(483) := b"1111111111111111_1111111111111111_1101101100111111_1100100101000000"; -- -0.14355795085430145
	pesos_i(484) := b"1111111111111111_1111111111111111_1101001000000110_1111101010000000"; -- -0.17958101630210876
	pesos_i(485) := b"0000000000000000_0000000000000000_0001100100110100_1111101110100000"; -- 0.09846470504999161
	pesos_i(486) := b"1111111111111111_1111111111111111_1001000111110000_0010010100000000"; -- -0.4299294352531433
	pesos_i(487) := b"0000000000000000_0000000000000000_0101110000010110_0100110110000000"; -- 0.3597153127193451
	pesos_i(488) := b"1111111111111111_1111111111111111_0000001111001111_0101110100000000"; -- -0.9851171374320984
	pesos_i(489) := b"1111111111111111_1111111111111111_1010110100011001_1011010010000000"; -- -0.32382652163505554
	pesos_i(490) := b"0000000000000000_0000000000000000_0010101111110001_1011100001000000"; -- 0.17165710031986237
	pesos_i(491) := b"0000000000000000_0000000000000000_0101011100011110_1100011110000000"; -- 0.3403134047985077
	pesos_i(492) := b"0000000000000000_0000000000000000_0110101000011100_1110000100000000"; -- 0.41450315713882446
	pesos_i(493) := b"1111111111111111_1111111111111111_1001101100110100_1001111100000000"; -- -0.3937283158302307
	pesos_i(494) := b"0000000000000000_0000000000000000_1001101110110111_0000011100000000"; -- 0.6082615256309509
	pesos_i(495) := b"1111111111111111_1111111111111111_1110101011000000_0010011010100000"; -- -0.08300551027059555
	pesos_i(496) := b"1111111111111111_1111111111111111_0110101101100101_1011000100000000"; -- -0.5804795622825623
	pesos_i(497) := b"0000000000000000_0000000000000000_0010100110010111_1111100010000000"; -- 0.16247513890266418
	pesos_i(498) := b"0000000000000000_0000000000000000_0110010011000110_1101100000000000"; -- 0.3936591148376465
	pesos_i(499) := b"1111111111111111_1111111111111111_0000111010001001_1000000100000000"; -- -0.9432143568992615
	pesos_i(500) := b"1111111111111111_1111111111111111_0000011010111111_1101100100000000"; -- -0.9736351370811462
	pesos_i(501) := b"0000000000000000_0000000000000000_0101000100010010_0000111100000000"; -- 0.31668180227279663
	pesos_i(502) := b"0000000000000000_0000000000000000_0000111111100101_1101101101010000"; -- 0.0621010847389698
	pesos_i(503) := b"0000000000000000_0000000000000000_0100100100111010_1010111010000000"; -- 0.2860516607761383
	pesos_i(504) := b"0000000000000000_0000000000000000_0111111110011111_0111110010000000"; -- 0.49852731823921204
	pesos_i(505) := b"0000000000000000_0000000000000000_1111100101101100_1111100100000000"; -- 0.9743190407752991
	pesos_i(506) := b"0000000000000000_0000000000000000_0011100000101011_1100001000000000"; -- 0.21941769123077393
	pesos_i(507) := b"1111111111111111_1111111111111111_0101111010001110_0001010000000000"; -- -0.6306445598602295
	pesos_i(508) := b"0000000000000000_0000000000000000_1000010010011111_1010101100000000"; -- 0.5180613398551941
	pesos_i(509) := b"1111111111111111_1111111111111111_0010011111010110_1001110100000000"; -- -0.8443815112113953
	pesos_i(510) := b"1111111111111111_1111111111111111_1100101101110100_0111011000000000"; -- -0.2052541971206665
	pesos_i(511) := b"0000000000000000_0000000000000000_0100001110010011_0000110010000000"; -- 0.2639625370502472
	pesos_i(512) := b"0000000000000000_0000000000000000_0101101100001011_1101011010000000"; -- 0.3556493818759918
	pesos_i(513) := b"1111111111111111_1111111111111111_0000110000101100_0001101100000000"; -- -0.9524520039558411
	pesos_i(514) := b"1111111111111111_1111111111111111_1111011001000100_1001011001110000"; -- -0.0380159355700016
	pesos_i(515) := b"1111111111111111_1111111111111111_1111110011010000_1001101110111000"; -- -0.012441890314221382
	pesos_i(516) := b"1111111111111111_1111111111111111_1010000101001000_0011000000000000"; -- -0.3699922561645508
	pesos_i(517) := b"0000000000000000_0000000000000000_1000111000011100_1001000100000000"; -- 0.5551233887672424
	pesos_i(518) := b"0000000000000000_0000000000000000_1010011000110100_0000100100000000"; -- 0.649231493473053
	pesos_i(519) := b"0000000000000000_0000000000000000_0101100100111100_1010001110000000"; -- 0.3485815227031708
	pesos_i(520) := b"1111111111111111_1111111111111111_0101010111110000_0111101100000000"; -- -0.6642993092536926
	pesos_i(521) := b"1111111111111111_1111111111111111_1000101111110111_1000100110000000"; -- -0.4532541334629059
	pesos_i(522) := b"1111111111111111_1111111111111111_1101100110111111_0001110011000000"; -- -0.1494276076555252
	pesos_i(523) := b"0000000000000000_0000000000000000_1001011011001110_0001100100000000"; -- 0.5890823006629944
	pesos_i(524) := b"0000000000000000_0000000000000000_0001010111100011_1010000110000000"; -- 0.08550462126731873
	pesos_i(525) := b"0000000000000000_0000000000000000_0011011011110110_1001101010000000"; -- 0.2147003710269928
	pesos_i(526) := b"0000000000000000_0000000000000000_0111000000111111_1110101000000000"; -- 0.43847525119781494
	pesos_i(527) := b"1111111111111111_1111111111111111_1101111110111000_0111110111000000"; -- -0.1260911375284195
	pesos_i(528) := b"0000000000000000_0000000000000000_0000001101000010_1100110010011100"; -- 0.01273802574723959
	pesos_i(529) := b"0000000000000000_0000000000000000_1001000110101111_0101101100000000"; -- 0.5690819621086121
	pesos_i(530) := b"0000000000000000_0000000000000000_0000011001101110_1011111101001000"; -- 0.025127368047833443
	pesos_i(531) := b"0000000000000000_0000000000000000_0101011101110000_0110001110000000"; -- 0.34155866503715515
	pesos_i(532) := b"0000000000000000_0000000000000000_0011100001101111_1000010110000000"; -- 0.22045168280601501
	pesos_i(533) := b"1111111111111111_1111111111111111_1110000110001110_1101000110000000"; -- -0.11891451478004456
	pesos_i(534) := b"1111111111111111_1111111111111111_1101011000011110_0000000110000000"; -- -0.16360464692115784
	pesos_i(535) := b"1111111111111111_1111111111111111_1110100100010001_1000101001100000"; -- -0.0895761027932167
	pesos_i(536) := b"1111111111111111_1111111111111111_1010110111101010_0100000110000000"; -- -0.3206442892551422
	pesos_i(537) := b"1111111111111111_1111111111111111_0101010110101000_1000110100000000"; -- -0.6653968691825867
	pesos_i(538) := b"0000000000000000_0000000000000000_0101001110100100_0011100010000000"; -- 0.3267245590686798
	pesos_i(539) := b"0000000000000000_0000000000000000_0010101010000110_0111100100000000"; -- 0.16611438989639282
	pesos_i(540) := b"0000000000000000_0000000000000000_1011000011111001_0011010100000000"; -- 0.6913025975227356
	pesos_i(541) := b"1111111111111111_1111111111111111_1101111011000100_0011001000000000"; -- -0.12981879711151123
	pesos_i(542) := b"1111111111111111_1111111111111111_0111010111101001_0111110000000000"; -- -0.5394060611724854
	pesos_i(543) := b"0000000000000000_0000000000000000_0000001100101111_1001111110011100"; -- 0.012445426546037197
	pesos_i(544) := b"0000000000000000_0000000000000000_1000000101011101_0001110100000000"; -- 0.505327045917511
	pesos_i(545) := b"1111111111111111_1111111111111111_0111110100000010_0101001000000000"; -- -0.5116833448410034
	pesos_i(546) := b"0000000000000000_0000000000000000_0100110000101110_1001111010000000"; -- 0.2975863516330719
	pesos_i(547) := b"1111111111111111_1111111111111111_1111000101110000_0010110110110000"; -- -0.056882042437791824
	pesos_i(548) := b"0000000000000000_0000000000000000_0100111000101011_1001111010000000"; -- 0.3053530752658844
	pesos_i(549) := b"0000000000000000_0000000000000000_1001100110000101_1110110100000000"; -- 0.5996997952461243
	pesos_i(550) := b"0000000000000000_0000000000000000_0000011101101000_1001010000110000"; -- 0.028939496725797653
	pesos_i(551) := b"1111111111111111_1111111111111111_1110010111101001_1010000110100000"; -- -0.10190381854772568
	pesos_i(552) := b"0000000000000000_0000000000000000_1000000110000111_0001000100000000"; -- 0.5059671998023987
	pesos_i(553) := b"0000000000000000_0000000000000000_1000100001011101_1101011000000000"; -- 0.5326818227767944
	pesos_i(554) := b"0000000000000000_0000000000000000_1010000011100011_0101100100000000"; -- 0.6284690499305725
	pesos_i(555) := b"0000000000000000_0000000000000000_0111111111101101_1010101100000000"; -- 0.4997202754020691
	pesos_i(556) := b"1111111111111111_1111111111111111_1000010000100110_1110111110000000"; -- -0.4837808907032013
	pesos_i(557) := b"1111111111111111_1111111111111111_1111111100110011_1111011011001011"; -- -0.003113341750577092
	pesos_i(558) := b"1111111111111111_1111111111111111_0110011100101110_1001110000000000"; -- -0.59694504737854
	pesos_i(559) := b"1111111111111111_1111111111111111_0110100000000011_0111010100000000"; -- -0.5936972498893738
	pesos_i(560) := b"0000000000000000_0000000000000000_0000011110101100_1100101111101000"; -- 0.029980415478348732
	pesos_i(561) := b"0000000000000000_0000000000000000_0010111110101001_1101001110000000"; -- 0.1861850917339325
	pesos_i(562) := b"1111111111111111_1111111111111111_0111011010011010_1001011000000000"; -- -0.5367037057876587
	pesos_i(563) := b"0000000000000000_0000000000000000_1000010000110110_1000001000000000"; -- 0.5164567232131958
	pesos_i(564) := b"1111111111111111_1111111111111111_0111000010111001_1000110100000000"; -- -0.5596687197685242
	pesos_i(565) := b"1111111111111111_1111111111111110_1110111010001111_0001110000000000"; -- -1.0681288242340088
	pesos_i(566) := b"0000000000000000_0000000000000000_0010010010111001_1110010011000000"; -- 0.14346151053905487
	pesos_i(567) := b"1111111111111111_1111111111111111_1001101011100001_1100101010000000"; -- -0.3949922025203705
	pesos_i(568) := b"1111111111111111_1111111111111111_0101101011001101_0011100000000000"; -- -0.6453061103820801
	pesos_i(569) := b"1111111111111111_1111111111111111_1100001110001000_0110111001000000"; -- -0.2361994832754135
	pesos_i(570) := b"1111111111111111_1111111111111111_1011100101010111_0010101010000000"; -- -0.27601370215415955
	pesos_i(571) := b"0000000000000000_0000000000000000_1111010011110110_1011000100000000"; -- 0.9568892121315002
	pesos_i(572) := b"1111111111111111_1111111111111111_1101100110110110_0110001100000000"; -- -0.14956074953079224
	pesos_i(573) := b"1111111111111111_1111111111111111_1101101010011110_0110100100000000"; -- -0.14602035284042358
	pesos_i(574) := b"0000000000000000_0000000000000000_0010101010110101_1110110100000000"; -- 0.16683846712112427
	pesos_i(575) := b"0000000000000000_0000000000000000_0111101001000010_1001111110000000"; -- 0.4775790870189667
	pesos_i(576) := b"1111111111111111_1111111111111111_1000001010101100_0000110010000000"; -- -0.4895622432231903
	pesos_i(577) := b"1111111111111111_1111111111111111_1100111111110110_0101011101000000"; -- -0.18764738738536835
	pesos_i(578) := b"0000000000000000_0000000000000000_0010011011111111_1110011101000000"; -- 0.1523422747850418
	pesos_i(579) := b"1111111111111111_1111111111111111_1110010100011111_1101000100000000"; -- -0.10498327016830444
	pesos_i(580) := b"1111111111111111_1111111111111111_1110101111011101_0100001000000000"; -- -0.07865512371063232
	pesos_i(581) := b"0000000000000000_0000000000000000_0111100111111001_1101101100000000"; -- 0.4764687418937683
	pesos_i(582) := b"1111111111111111_1111111111111111_0101010101011100_0110111100000000"; -- -0.6665583252906799
	pesos_i(583) := b"1111111111111111_1111111111111111_0111101110010010_1011001000000000"; -- -0.517292857170105
	pesos_i(584) := b"1111111111111111_1111111111111111_1010010001101001_1010111110000000"; -- -0.3577623665332794
	pesos_i(585) := b"1111111111111111_1111111111111111_0111001110111000_1111001100000000"; -- -0.5479591488838196
	pesos_i(586) := b"0000000000000000_0000000000000000_0010011010000111_1001111001000000"; -- 0.1505068689584732
	pesos_i(587) := b"0000000000000000_0000000000000000_0111111100111110_1110010010000000"; -- 0.4970534145832062
	pesos_i(588) := b"1111111111111111_1111111111111111_1000000101111111_1000111100000000"; -- -0.4941473603248596
	pesos_i(589) := b"1111111111111111_1111111111111111_1011010010111111_0100111110000000"; -- -0.29395583271980286
	pesos_i(590) := b"1111111111111111_1111111111111111_1111010011111111_0000100100000000"; -- -0.04298347234725952
	pesos_i(591) := b"1111111111111111_1111111111111111_1110011111111101_1100000001100000"; -- -0.09378430992364883
	pesos_i(592) := b"1111111111111111_1111111111111111_1011011010000011_1110110110000000"; -- -0.28704944252967834
	pesos_i(593) := b"0000000000000000_0000000000000001_0000011111110101_1100100000000000"; -- 1.0310940742492676
	pesos_i(594) := b"1111111111111111_1111111111111111_1111110101111101_0111010111111000"; -- -0.009804369881749153
	pesos_i(595) := b"1111111111111111_1111111111111111_1111100001000111_0111100101111000"; -- -0.03015938587486744
	pesos_i(596) := b"1111111111111111_1111111111111111_0100110111100000_1010110000000000"; -- -0.6957905292510986
	pesos_i(597) := b"1111111111111111_1111111111111111_0110000000111000_1111111100000000"; -- -0.6241303086280823
	pesos_i(598) := b"1111111111111111_1111111111111111_1011000111100110_0000000000000000"; -- -0.305084228515625
	pesos_i(599) := b"1111111111111111_1111111111111111_0111011010111110_1000000000000000"; -- -0.5361557006835938
	pesos_i(600) := b"1111111111111111_1111111111111111_1000101111010011_0011000110000000"; -- -0.4538086950778961
	pesos_i(601) := b"0000000000000000_0000000000000000_0000010010100011_0110001101010000"; -- 0.018118102103471756
	pesos_i(602) := b"1111111111111111_1111111111111111_0010100110001010_1000000100000000"; -- -0.837730348110199
	pesos_i(603) := b"1111111111111111_1111111111111111_1011110101000101_1000000110000000"; -- -0.2606581747531891
	pesos_i(604) := b"0000000000000000_0000000000000000_0000011111010110_1110010110100000"; -- 0.03062281757593155
	pesos_i(605) := b"1111111111111111_1111111111111111_0011111011000111_1101110000000000"; -- -0.7547628879547119
	pesos_i(606) := b"0000000000000000_0000000000000000_0110100100101001_0011101000000000"; -- 0.4107853174209595
	pesos_i(607) := b"0000000000000000_0000000000000000_0110010010110100_0000010100000000"; -- 0.3933718800544739
	pesos_i(608) := b"1111111111111111_1111111111111111_1111010110111100_0110010000000000"; -- -0.04009413719177246
	pesos_i(609) := b"0000000000000000_0000000000000000_0000101101110010_0100011101000000"; -- 0.04471249878406525
	pesos_i(610) := b"0000000000000000_0000000000000000_0011000111011100_0001001101000000"; -- 0.19476433098316193
	pesos_i(611) := b"1111111111111111_1111111111111111_1111100110001001_0010000101000000"; -- -0.025251314043998718
	pesos_i(612) := b"1111111111111111_1111111111111111_1000011000011100_1011111110000000"; -- -0.4761238396167755
	pesos_i(613) := b"1111111111111111_1111111111111111_1011001001101011_0010101110000000"; -- -0.30305221676826477
	pesos_i(614) := b"1111111111111111_1111111111111111_1111001001011101_0110110001100000"; -- -0.05326197296380997
	pesos_i(615) := b"0000000000000000_0000000000000000_0111000001100100_1001011100000000"; -- 0.4390348792076111
	pesos_i(616) := b"1111111111111111_1111111111111111_0110011111011110_0000001000000000"; -- -0.5942686796188354
	pesos_i(617) := b"0000000000000000_0000000000000000_0000000101010010_1100110111101100"; -- 0.005169744603335857
	pesos_i(618) := b"1111111111111111_1111111111111111_1111111111101110_0101010010101110"; -- -0.0002696109004318714
	pesos_i(619) := b"1111111111111111_1111111111111111_1100100010100110_0001100000000000"; -- -0.2162156105041504
	pesos_i(620) := b"0000000000000000_0000000000000000_1011110110111000_1110101100000000"; -- 0.7411028742790222
	pesos_i(621) := b"0000000000000000_0000000000000000_0011110110100110_1000110011000000"; -- 0.24082259833812714
	pesos_i(622) := b"0000000000000000_0000000000000000_0111011111100010_1111010100000000"; -- 0.46830683946609497
	pesos_i(623) := b"1111111111111111_1111111111111111_0100111000010001_1110000100000000"; -- -0.695039689540863
	pesos_i(624) := b"1111111111111111_1111111111111111_0011101101111001_1100110000000000"; -- -0.7676727771759033
	pesos_i(625) := b"0000000000000000_0000000000000000_0100010100010110_0000010100000000"; -- 0.2698672413825989
	pesos_i(626) := b"0000000000000000_0000000000000000_0011101000101000_0001011100000000"; -- 0.22717422246932983
	pesos_i(627) := b"1111111111111111_1111111111111111_1000111010011001_0010110010000000"; -- -0.442975252866745
	pesos_i(628) := b"1111111111111111_1111111111111111_0001010100010010_1010001100000000"; -- -0.9176843762397766
	pesos_i(629) := b"0000000000000000_0000000000000000_0101001011101000_0000001110000000"; -- 0.3238527476787567
	pesos_i(630) := b"1111111111111111_1111111111111111_1110010100101101_1001010011000000"; -- -0.10477323830127716
	pesos_i(631) := b"0000000000000000_0000000000000000_0011101010100001_0001111000000000"; -- 0.22902095317840576
	pesos_i(632) := b"0000000000000000_0000000000000000_0111011111110001_1001000000000000"; -- 0.46852970123291016
	pesos_i(633) := b"0000000000000000_0000000000000000_1010101101110011_0101110000000000"; -- 0.6697289943695068
	pesos_i(634) := b"0000000000000000_0000000000000000_0010001010111101_1110010100000000"; -- 0.13571006059646606
	pesos_i(635) := b"1111111111111111_1111111111111111_1010100100101010_1110010100000000"; -- -0.33918923139572144
	pesos_i(636) := b"0000000000000000_0000000000000000_1000010000100110_1110101000000000"; -- 0.5162187814712524
	pesos_i(637) := b"1111111111111111_1111111111111111_0111110010110010_0011010100000000"; -- -0.5129057765007019
	pesos_i(638) := b"1111111111111111_1111111111111111_1001010010010000_0000111100000000"; -- -0.41967684030532837
	pesos_i(639) := b"1111111111111111_1111111111111111_1110000010110101_1100111000100000"; -- -0.12222587317228317
	pesos_i(640) := b"0000000000000000_0000000000000000_1000110101001110_1000100000000000"; -- 0.5519795417785645
	pesos_i(641) := b"1111111111111111_1111111111111111_1111100110110001_1000110010011000"; -- -0.02463456429541111
	pesos_i(642) := b"1111111111111111_1111111111111111_1000110101111111_0010110000000000"; -- -0.4472782611846924
	pesos_i(643) := b"0000000000000000_0000000000000000_1000001001100001_0110010000000000"; -- 0.50929856300354
	pesos_i(644) := b"1111111111111111_1111111111111111_1011111001110110_0011011000000000"; -- -0.25600874423980713
	pesos_i(645) := b"1111111111111111_1111111111111111_1100011010101110_1100001000000000"; -- -0.22389590740203857
	pesos_i(646) := b"0000000000000000_0000000000000000_1000110001100001_0111001100000000"; -- 0.5483619570732117
	pesos_i(647) := b"0000000000000000_0000000000000000_0110110011101011_1000111100000000"; -- 0.4254693388938904
	pesos_i(648) := b"1111111111111111_1111111111111111_0101111101110010_1000011100000000"; -- -0.6271587014198303
	pesos_i(649) := b"1111111111111111_1111111111111111_0111100000001111_0001101100000000"; -- -0.5310195088386536
	pesos_i(650) := b"0000000000000000_0000000000000000_0101011111100101_0000010000000000"; -- 0.3433382511138916
	pesos_i(651) := b"0000000000000000_0000000000000000_0000110011110001_1001111100110000"; -- 0.05056185647845268
	pesos_i(652) := b"0000000000000000_0000000000000000_0100110100000000_1100111110000000"; -- 0.3007936179637909
	pesos_i(653) := b"0000000000000000_0000000000000000_0100111111011000_1000010110000000"; -- 0.3118976056575775
	pesos_i(654) := b"0000000000000000_0000000000000000_0001010001110011_1000001100000000"; -- 0.07988756895065308
	pesos_i(655) := b"1111111111111111_1111111111111111_1100011001010001_0100101010000000"; -- -0.22532209753990173
	pesos_i(656) := b"0000000000000000_0000000000000000_0110011100011101_0111001100000000"; -- 0.40279310941696167
	pesos_i(657) := b"0000000000000000_0000000000000000_0100111100110000_1000100100000000"; -- 0.30933433771133423
	pesos_i(658) := b"1111111111111111_1111111111111111_1010110010010000_0101011000000000"; -- -0.3259226083755493
	pesos_i(659) := b"1111111111111111_1111111111111111_1111110111110110_1100001000011100"; -- -0.007953518070280552
	pesos_i(660) := b"0000000000000000_0000000000000000_0110001001100111_0100100110000000"; -- 0.3843885362148285
	pesos_i(661) := b"1111111111111111_1111111111111111_0111011101110111_0100111100000000"; -- -0.5333357453346252
	pesos_i(662) := b"1111111111111111_1111111111111111_0111011101100101_0000110100000000"; -- -0.5336143374443054
	pesos_i(663) := b"0000000000000000_0000000000000000_0001010101001000_0110010111100000"; -- 0.08313595503568649
	pesos_i(664) := b"1111111111111111_1111111111111111_1011010001111010_1101111000000000"; -- -0.29500019550323486
	pesos_i(665) := b"1111111111111111_1111111111111111_1000100100100101_0001001000000000"; -- -0.46427810192108154
	pesos_i(666) := b"1111111111111111_1111111111111111_1010010000111101_1010011010000000"; -- -0.3584342896938324
	pesos_i(667) := b"0000000000000000_0000000000000000_0000011100111001_0000000000111000"; -- 0.028213514015078545
	pesos_i(668) := b"0000000000000000_0000000000000000_0001100111100110_0110000001000000"; -- 0.10117150843143463
	pesos_i(669) := b"0000000000000000_0000000000000000_0101010111101001_1100101100000000"; -- 0.3355986475944519
	pesos_i(670) := b"1111111111111111_1111111111111111_0101101100110100_1001100100000000"; -- -0.6437286734580994
	pesos_i(671) := b"1111111111111111_1111111111111111_1111100101001101_0110101110111000"; -- -0.0261624027043581
	pesos_i(672) := b"0000000000000000_0000000000000000_0011101010001011_1011110101000000"; -- 0.22869475185871124
	pesos_i(673) := b"1111111111111111_1111111111111111_1110011010011101_1000011011100000"; -- -0.09915883094072342
	pesos_i(674) := b"0000000000000000_0000000000000000_1000110011101111_1110111000000000"; -- 0.550536036491394
	pesos_i(675) := b"0000000000000000_0000000000000000_1000000010110110_0001110100000000"; -- 0.5027788281440735
	pesos_i(676) := b"0000000000000000_0000000000000000_1010000111101100_0000010100000000"; -- 0.6325076222419739
	pesos_i(677) := b"0000000000000000_0000000000000000_1001100101000011_0100001100000000"; -- 0.5986825823783875
	pesos_i(678) := b"0000000000000000_0000000000000000_0010101111101110_0101110010000000"; -- 0.17160585522651672
	pesos_i(679) := b"0000000000000000_0000000000000000_0011011101011100_1100011000000000"; -- 0.21625936031341553
	pesos_i(680) := b"0000000000000000_0000000000000000_1110101000011110_0101111100000000"; -- 0.9145259261131287
	pesos_i(681) := b"0000000000000000_0000000000000000_0111011100101010_1010000110000000"; -- 0.4654942452907562
	pesos_i(682) := b"0000000000000000_0000000000000000_0100110111101011_0101010010000000"; -- 0.304372102022171
	pesos_i(683) := b"0000000000000000_0000000000000000_0011111010011011_0111101001000000"; -- 0.2445598989725113
	pesos_i(684) := b"1111111111111111_1111111111111111_0011001111000000_0100101100000000"; -- -0.7978470921516418
	pesos_i(685) := b"0000000000000000_0000000000000000_0011000101011001_0101011110000000"; -- 0.19276949763298035
	pesos_i(686) := b"0000000000000000_0000000000000000_0000101001010100_0010001110100000"; -- 0.04034636169672012
	pesos_i(687) := b"1111111111111111_1111111111111111_1010111011000111_1001110000000000"; -- -0.31726670265197754
	pesos_i(688) := b"1111111111111111_1111111111111111_1011110000111111_0101111000000000"; -- -0.2646580934524536
	pesos_i(689) := b"0000000000000000_0000000000000000_0001110110011100_0101001111100000"; -- 0.11566662043333054
	pesos_i(690) := b"1111111111111111_1111111111111111_1110000001111000_0101111000100000"; -- -0.12316333502531052
	pesos_i(691) := b"0000000000000000_0000000000000000_1100101100100010_0000010000000000"; -- 0.7934877872467041
	pesos_i(692) := b"1111111111111111_1111111111111111_1111000111010101_0000110101100000"; -- -0.05534283071756363
	pesos_i(693) := b"1111111111111111_1111111111111111_0101101011100100_1000001100000000"; -- -0.6449506878852844
	pesos_i(694) := b"1111111111111111_1111111111111111_1111111001100101_1001011000001100"; -- -0.0062624188140034676
	pesos_i(695) := b"1111111111111111_1111111111111111_1000000101011011_1101100010000000"; -- -0.49469229578971863
	pesos_i(696) := b"1111111111111111_1111111111111111_1001111111011110_1111111100000000"; -- -0.3755035996437073
	pesos_i(697) := b"1111111111111111_1111111111111111_1010010010001110_0010000110000000"; -- -0.357206255197525
	pesos_i(698) := b"0000000000000000_0000000000000000_0000111111011010_0100010011000000"; -- 0.06192426383495331
	pesos_i(699) := b"0000000000000000_0000000000000000_0111010101100000_1000000010000000"; -- 0.45850375294685364
	pesos_i(700) := b"1111111111111111_1111111111111111_0111110111000001_1011111000000000"; -- -0.5087624788284302
	pesos_i(701) := b"1111111111111111_1111111111111111_1111001010010101_1101010110110000"; -- -0.05240120366215706
	pesos_i(702) := b"0000000000000000_0000000000000000_0100100101100011_1110100000000000"; -- 0.2866806983947754
	pesos_i(703) := b"0000000000000000_0000000000000000_1001100101110110_0101001100000000"; -- 0.5994617342948914
	pesos_i(704) := b"0000000000000000_0000000000000000_0011011101111000_1001010111000000"; -- 0.21668373048305511
	pesos_i(705) := b"0000000000000000_0000000000000000_0000011101011000_1101110101000000"; -- 0.028699710965156555
	pesos_i(706) := b"1111111111111111_1111111111111111_1111001010111000_1011110010000000"; -- -0.05186864733695984
	pesos_i(707) := b"1111111111111111_1111111111111111_1100100010010001_1110011101000000"; -- -0.2165236920118332
	pesos_i(708) := b"0000000000000000_0000000000000000_0000010010000110_1000110100100000"; -- 0.017678089439868927
	pesos_i(709) := b"0000000000000000_0000000000000000_0000011110101011_0101001100110000"; -- 0.029957961291074753
	pesos_i(710) := b"1111111111111111_1111111111111111_1010011101110000_1110010110000000"; -- -0.34593358635902405
	pesos_i(711) := b"1111111111111111_1111111111111111_1001001011000010_1011110000000000"; -- -0.4267160892486572
	pesos_i(712) := b"1111111111111111_1111111111111111_1001111001001010_0110111100000000"; -- -0.38167673349380493
	pesos_i(713) := b"1111111111111111_1111111111111111_1100100110011010_1101010001000000"; -- -0.21248124539852142
	pesos_i(714) := b"0000000000000000_0000000000000000_0010110000101010_1100111001000000"; -- 0.17252816259860992
	pesos_i(715) := b"0000000000000000_0000000000000000_1000100100111011_0000111100000000"; -- 0.5360574126243591
	pesos_i(716) := b"1111111111111111_1111111111111111_0111011101101010_0100110000000000"; -- -0.5335342884063721
	pesos_i(717) := b"1111111111111111_1111111111111111_1010111001110011_0001101000000000"; -- -0.31855618953704834
	pesos_i(718) := b"1111111111111111_1111111111111111_1110000100101101_1111000001000000"; -- -0.12039278447628021
	pesos_i(719) := b"0000000000000000_0000000000000000_0001111100111000_0001100000000000"; -- 0.12194967269897461
	pesos_i(720) := b"1111111111111111_1111111111111111_1100010101011100_1011010110000000"; -- -0.22905412316322327
	pesos_i(721) := b"0000000000000000_0000000000000001_0001001110111011_1111000000000000"; -- 1.0770864486694336
	pesos_i(722) := b"0000000000000000_0000000000000000_0001001101111011_0001110011100000"; -- 0.07609730213880539
	pesos_i(723) := b"0000000000000000_0000000000000000_0011110111110101_1000010000000000"; -- 0.24202752113342285
	pesos_i(724) := b"0000000000000000_0000000000000000_0010111001111000_0111001100000000"; -- 0.18152540922164917
	pesos_i(725) := b"1111111111111111_1111111111111111_1101110111000000_0100001011000000"; -- -0.13378508388996124
	pesos_i(726) := b"1111111111111111_1111111111111111_1000011100011001_1110101100000000"; -- -0.4722607731819153
	pesos_i(727) := b"1111111111111111_1111111111111111_0101101110001011_1010110100000000"; -- -0.6423999667167664
	pesos_i(728) := b"1111111111111111_1111111111111111_1000101111111101_0111101110000000"; -- -0.45316341519355774
	pesos_i(729) := b"0000000000000000_0000000000000000_1001110100001111_1001111000000000"; -- 0.613519549369812
	pesos_i(730) := b"1111111111111111_1111111111111111_0100001101110000_0110000000000000"; -- -0.7365665435791016
	pesos_i(731) := b"1111111111111111_1111111111111111_0101010110011011_1011101000000000"; -- -0.6655925512313843
	pesos_i(732) := b"0000000000000000_0000000000000000_0010010111110010_0000101101000000"; -- 0.14822454750537872
	pesos_i(733) := b"1111111111111111_1111111111111111_0110111101011001_0110000100000000"; -- -0.5650424361228943
	pesos_i(734) := b"0000000000000000_0000000000000000_0101100001111100_0011111010000000"; -- 0.34564581513404846
	pesos_i(735) := b"1111111111111111_1111111111111111_1000010110100010_1100000100000000"; -- -0.47798532247543335
	pesos_i(736) := b"1111111111111111_1111111111111111_1011111001101100_0110001100000000"; -- -0.25615864992141724
	pesos_i(737) := b"1111111111111111_1111111111111111_1101001110011100_1100101010000000"; -- -0.17338880896568298
	pesos_i(738) := b"1111111111111111_1111111111111111_1110010000111110_1011010000100000"; -- -0.10841821879148483
	pesos_i(739) := b"0000000000000000_0000000000000000_0100010101111111_1111101100000000"; -- 0.2714840769767761
	pesos_i(740) := b"1111111111111111_1111111111111111_0111111001000100_0100001000000000"; -- -0.5067709684371948
	pesos_i(741) := b"1111111111111111_1111111111111111_1001111110010111_1110011010000000"; -- -0.3765884339809418
	pesos_i(742) := b"0000000000000000_0000000000000000_0000011100111100_0100001101111000"; -- 0.02826329879462719
	pesos_i(743) := b"1111111111111111_1111111111111111_1101010111011001_1110011010000000"; -- -0.16464385390281677
	pesos_i(744) := b"0000000000000000_0000000000000000_0010000011100010_0001111101000000"; -- 0.12845034897327423
	pesos_i(745) := b"0000000000000000_0000000000000000_0010100011101110_1000110001000000"; -- 0.15988995134830475
	pesos_i(746) := b"0000000000000000_0000000000000000_0010011110011111_1011111010000000"; -- 0.1547812521457672
	pesos_i(747) := b"1111111111111111_1111111111111111_1011010000111000_0100111100000000"; -- -0.29601579904556274
	pesos_i(748) := b"0000000000000000_0000000000000000_1011010101010101_1101000100000000"; -- 0.7083407044410706
	pesos_i(749) := b"0000000000000000_0000000000000000_0111101001011111_0011011110000000"; -- 0.47801539301872253
	pesos_i(750) := b"1111111111111111_1111111111111111_1011000011110110_1101100100000000"; -- -0.30873340368270874
	pesos_i(751) := b"1111111111111111_1111111111111111_0011000101000100_0010111000000000"; -- -0.8075534105300903
	pesos_i(752) := b"1111111111111111_1111111111111111_1000101100011101_1000011010000000"; -- -0.4565807282924652
	pesos_i(753) := b"1111111111111111_1111111111111111_1001110010100111_0010011110000000"; -- -0.38807442784309387
	pesos_i(754) := b"0000000000000000_0000000000000000_1001111011100110_0000001000000000"; -- 0.6206971406936646
	pesos_i(755) := b"1111111111111111_1111111111111111_1011100011110011_0011111110000000"; -- -0.27753832936286926
	pesos_i(756) := b"1111111111111111_1111111111111111_0100101011011001_1111011100000000"; -- -0.707611620426178
	pesos_i(757) := b"0000000000000000_0000000000000000_0101001011010100_1101110010000000"; -- 0.323560506105423
	pesos_i(758) := b"1111111111111111_1111111111111111_1111110001001011_0111111111000100"; -- -0.01447297539561987
	pesos_i(759) := b"1111111111111111_1111111111111111_1000000000101011_1010011110000000"; -- -0.4993338882923126
	pesos_i(760) := b"0000000000000000_0000000000000000_0011111111110111_1111100011000000"; -- 0.24987749755382538
	pesos_i(761) := b"0000000000000000_0000000000000000_0111001001110111_0010110110000000"; -- 0.4471310079097748
	pesos_i(762) := b"0000000000000000_0000000000000000_0001011001010001_0011101010100000"; -- 0.08717695623636246
	pesos_i(763) := b"1111111111111111_1111111111111111_1111101001101010_0100011011000000"; -- -0.02181585133075714
	pesos_i(764) := b"0000000000000000_0000000000000000_0111010101101110_1001110110000000"; -- 0.4587191045284271
	pesos_i(765) := b"1111111111111111_1111111111111111_1001011011100110_0110000000000000"; -- -0.41054725646972656
	pesos_i(766) := b"1111111111111111_1111111111111111_1111001001101001_0100000110110000"; -- -0.053081411868333817
	pesos_i(767) := b"1111111111111111_1111111111111111_1001101101010100_1000011010000000"; -- -0.3932414948940277
	pesos_i(768) := b"0000000000000000_0000000000000000_0001011101110011_0101010011000000"; -- 0.09160356223583221
	pesos_i(769) := b"1111111111111111_1111111111111111_1111000001111010_0011111011100000"; -- -0.06063468009233475
	pesos_i(770) := b"1111111111111111_1111111111111111_1111011001101001_0001100111100000"; -- -0.03745878487825394
	pesos_i(771) := b"0000000000000000_0000000000000000_0011110110101101_0101101100000000"; -- 0.24092644453048706
	pesos_i(772) := b"1111111111111111_1111111111111111_1101001011010000_0110001001000000"; -- -0.17650781571865082
	pesos_i(773) := b"1111111111111111_1111111111111111_1010001110011001_0101001000000000"; -- -0.3609417676925659
	pesos_i(774) := b"0000000000000000_0000000000000000_0101000000100001_0110111100000000"; -- 0.31301015615463257
	pesos_i(775) := b"0000000000000000_0000000000000000_0011001100100000_1010100000000000"; -- 0.19971704483032227
	pesos_i(776) := b"1111111111111111_1111111111111111_1100000101010001_0100100111000000"; -- -0.24485339224338531
	pesos_i(777) := b"1111111111111111_1111111111111111_1111000001111000_0111010100010000"; -- -0.06066196784377098
	pesos_i(778) := b"1111111111111111_1111111111111111_1111111010100001_1111101100001000"; -- -0.005340872332453728
	pesos_i(779) := b"1111111111111111_1111111111111111_1100001010100101_0011111101000000"; -- -0.23966602981090546
	pesos_i(780) := b"0000000000000000_0000000000000000_0100011110010000_0000000110000000"; -- 0.27954110503196716
	pesos_i(781) := b"0000000000000000_0000000000000000_0010011100001010_1101101110000000"; -- 0.1525094211101532
	pesos_i(782) := b"0000000000000000_0000000000000000_0000001100110011_1100110001010100"; -- 0.012509127147495747
	pesos_i(783) := b"1111111111111111_1111111111111111_1010101001000110_1011001100000000"; -- -0.3348587155342102
	pesos_i(784) := b"0000000000000000_0000000000000000_0000001010100100_0010000010010100"; -- 0.010316883213818073
	pesos_i(785) := b"0000000000000000_0000000000000000_0100000100011001_0111111000000000"; -- 0.2542952299118042
	pesos_i(786) := b"1111111111111111_1111111111111111_1101011001010101_1001000111000000"; -- -0.1627568155527115
	pesos_i(787) := b"1111111111111111_1111111111111111_1111101001010011_1101011000110000"; -- -0.02215825393795967
	pesos_i(788) := b"0000000000000000_0000000000000000_0011000010000001_1010000010000000"; -- 0.18947795033454895
	pesos_i(789) := b"1111111111111111_1111111111111111_0111100010011001_1001010000000000"; -- -0.5289065837860107
	pesos_i(790) := b"1111111111111111_1111111111111111_1110011001010110_0001001101000000"; -- -0.10024909675121307
	pesos_i(791) := b"1111111111111111_1111111111111111_1101110111101001_1111100100000000"; -- -0.13314861059188843
	pesos_i(792) := b"1111111111111111_1111111111111111_1001101101010110_0111110000000000"; -- -0.39321160316467285
	pesos_i(793) := b"1111111111111111_1111111111111111_1100010101000000_0100101011000000"; -- -0.22948773205280304
	pesos_i(794) := b"1111111111111111_1111111111111111_1101110010001011_1010011011000000"; -- -0.1384940892457962
	pesos_i(795) := b"1111111111111111_1111111111111111_1110001100011000_0100001000000000"; -- -0.11291110515594482
	pesos_i(796) := b"1111111111111111_1111111111111111_1111010000100011_1000001100000000"; -- -0.046333134174346924
	pesos_i(797) := b"0000000000000000_0000000000000000_0010100000100000_0110011110000000"; -- 0.15674445033073425
	pesos_i(798) := b"1111111111111111_1111111111111111_1101001110001011_0000111101000000"; -- -0.17365936934947968
	pesos_i(799) := b"0000000000000000_0000000000000000_0011010000100100_0101001001000000"; -- 0.20367921888828278
	pesos_i(800) := b"0000000000000000_0000000000000000_0010101001010101_1101000000000000"; -- 0.16537189483642578
	pesos_i(801) := b"0000000000000000_0000000000000000_0000101000110101_1010101101010000"; -- 0.039881426841020584
	pesos_i(802) := b"0000000000000000_0000000000000000_0110001101000101_1111111110000000"; -- 0.3877868354320526
	pesos_i(803) := b"0000000000000000_0000000000000000_0101001000010101_1010110000000000"; -- 0.32064318656921387
	pesos_i(804) := b"0000000000000000_0000000000000000_0111010110011011_1100111100000000"; -- 0.459408700466156
	pesos_i(805) := b"0000000000000000_0000000000000000_0000100111100100_1111101111100000"; -- 0.0386502668261528
	pesos_i(806) := b"0000000000000000_0000000000000000_0010000001000000_0011001111000000"; -- 0.12597964704036713
	pesos_i(807) := b"0000000000000000_0000000000000000_0011001000101100_1000100000000000"; -- 0.19599199295043945
	pesos_i(808) := b"0000000000000000_0000000000000000_1000000000111110_0101111000000000"; -- 0.5009516477584839
	pesos_i(809) := b"0000000000000000_0000000000000000_0010101000000111_1110001100000000"; -- 0.1641828417778015
	pesos_i(810) := b"1111111111111111_1111111111111111_1111111100110010_0100111100010100"; -- -0.003138597123324871
	pesos_i(811) := b"0000000000000000_0000000000000000_0010001100011010_0100011111000000"; -- 0.13711975514888763
	pesos_i(812) := b"1111111111111111_1111111111111111_1010011110000111_0111101010000000"; -- -0.3455890119075775
	pesos_i(813) := b"0000000000000000_0000000000000000_0011110100110111_0001100101000000"; -- 0.23912198841571808
	pesos_i(814) := b"0000000000000000_0000000000000000_0010110110010000_0010110101000000"; -- 0.1779812127351761
	pesos_i(815) := b"1111111111111111_1111111111111111_1111100110011011_1100100100111000"; -- -0.024966644123196602
	pesos_i(816) := b"1111111111111111_1111111111111111_1110011101110110_0011110001000000"; -- -0.09585212171077728
	pesos_i(817) := b"1111111111111111_1111111111111111_1110001000100001_0101001001000000"; -- -0.11667905747890472
	pesos_i(818) := b"1111111111111111_1111111111111111_1110001111001000_1101011101100000"; -- -0.1102166548371315
	pesos_i(819) := b"0000000000000000_0000000000000000_0001001010101101_0111111010100000"; -- 0.07295981794595718
	pesos_i(820) := b"0000000000000000_0000000000000000_0011100100110111_0010001110000000"; -- 0.22349759936332703
	pesos_i(821) := b"1111111111111111_1111111111111111_1001000111101010_1000011010000000"; -- -0.4300151765346527
	pesos_i(822) := b"0000000000000000_0000000000000000_0010101011000111_1111001001000000"; -- 0.16711343824863434
	pesos_i(823) := b"1111111111111111_1111111111111111_1111101000110110_0010000001000000"; -- -0.022611603140830994
	pesos_i(824) := b"1111111111111111_1111111111111111_1101100000101101_1000000110000000"; -- -0.1555556356906891
	pesos_i(825) := b"0000000000000000_0000000000000000_0000010010100111_1101100110111000"; -- 0.018186194822192192
	pesos_i(826) := b"0000000000000000_0000000000000000_0000100101010100_1100011010110000"; -- 0.03644983097910881
	pesos_i(827) := b"0000000000000000_0000000000000000_0001110000111000_0001101010000000"; -- 0.11023107171058655
	pesos_i(828) := b"1111111111111111_1111111111111111_1010000010011010_0110001010000000"; -- -0.3726442754268646
	pesos_i(829) := b"0000000000000000_0000000000000000_0011010111101001_1001011101000000"; -- 0.21059556305408478
	pesos_i(830) := b"1111111111111111_1111111111111111_1101111110101001_1000110000000000"; -- -0.12631916999816895
	pesos_i(831) := b"0000000000000000_0000000000000000_0011110111111110_1111011010000000"; -- 0.24217167496681213
	pesos_i(832) := b"1111111111111111_1111111111111111_1110011001011000_1101000110100000"; -- -0.10020723193883896
	pesos_i(833) := b"0000000000000000_0000000000000000_0001011001101001_0010110101100000"; -- 0.08754237741231918
	pesos_i(834) := b"0000000000000000_0000000000000000_0000001110101110_1110111100111100"; -- 0.014388038776814938
	pesos_i(835) := b"0000000000000000_0000000000000000_0010000101111110_0010110011000000"; -- 0.1308315247297287
	pesos_i(836) := b"1111111111111111_1111111111111111_1010100010111010_1110110000000000"; -- -0.340897798538208
	pesos_i(837) := b"1111111111111111_1111111111111111_1111111100111000_1011100010010100"; -- -0.0030407560989260674
	pesos_i(838) := b"1111111111111111_1111111111111111_1110101010111000_0010110000000000"; -- -0.08312726020812988
	pesos_i(839) := b"1111111111111111_1111111111111111_1001011000010011_1110010110000000"; -- -0.41375890374183655
	pesos_i(840) := b"1111111111111111_1111111111111111_1011010100011110_1001010100000000"; -- -0.29250210523605347
	pesos_i(841) := b"1111111111111111_1111111111111111_1110101111001001_1010010111100000"; -- -0.07895434647798538
	pesos_i(842) := b"0000000000000000_0000000000000000_0010100111110000_0011110101000000"; -- 0.1638220101594925
	pesos_i(843) := b"0000000000000000_0000000000000000_0100100001101001_1010010100000000"; -- 0.28286200761795044
	pesos_i(844) := b"1111111111111111_1111111111111111_1110010001001010_1001100001000000"; -- -0.10823677480220795
	pesos_i(845) := b"1111111111111111_1111111111111111_1101000010000101_1001100100000000"; -- -0.18546146154403687
	pesos_i(846) := b"0000000000000000_0000000000000000_0000100101101000_1001001101000000"; -- 0.036751940846443176
	pesos_i(847) := b"0000000000000000_0000000000000000_0001000000000000_0100100110100000"; -- 0.06250438839197159
	pesos_i(848) := b"0000000000000000_0000000000000000_0000011011101101_1101100100100000"; -- 0.027066774666309357
	pesos_i(849) := b"0000000000000000_0000000000000000_0111010010101001_1101000000000000"; -- 0.4557161331176758
	pesos_i(850) := b"1111111111111111_1111111111111111_1111100010011100_1011111111111000"; -- -0.028858186677098274
	pesos_i(851) := b"0000000000000000_0000000000000000_0011010111110111_0011100000000000"; -- 0.21080350875854492
	pesos_i(852) := b"0000000000000000_0000000000000000_0000100000111101_0110010101110000"; -- 0.032186832278966904
	pesos_i(853) := b"0000000000000000_0000000000000000_0000000100000000_1100000001111100"; -- 0.003917722962796688
	pesos_i(854) := b"1111111111111111_1111111111111111_1011110100000110_0000000110000000"; -- -0.26162710785865784
	pesos_i(855) := b"1111111111111111_1111111111111111_1110000110111110_0001111101100000"; -- -0.11819270998239517
	pesos_i(856) := b"1111111111111111_1111111111111111_1111001010001011_1011011101100000"; -- -0.05255559831857681
	pesos_i(857) := b"0000000000000000_0000000000000000_0101101001010000_0100110110000000"; -- 0.3527878224849701
	pesos_i(858) := b"1111111111111111_1111111111111111_1001100011100101_1111101110000000"; -- -0.4027407467365265
	pesos_i(859) := b"1111111111111111_1111111111111111_1100101111011100_1010001000000000"; -- -0.2036646604537964
	pesos_i(860) := b"0000000000000000_0000000000000000_0011000010110000_0010000001000000"; -- 0.190187469124794
	pesos_i(861) := b"1111111111111111_1111111111111111_1011110011101111_1111100100000000"; -- -0.2619633078575134
	pesos_i(862) := b"0000000000000000_0000000000000000_0100101011011010_1011100000000000"; -- 0.29239988327026367
	pesos_i(863) := b"1111111111111111_1111111111111111_1010011110000010_0110101000000000"; -- -0.3456662893295288
	pesos_i(864) := b"1111111111111111_1111111111111111_1100111011001000_1010010111000000"; -- -0.19225086271762848
	pesos_i(865) := b"0000000000000000_0000000000000000_0010110101001001_0101101000000000"; -- 0.17690050601959229
	pesos_i(866) := b"1111111111111111_1111111111111111_1110000101001110_0100100000100000"; -- -0.11989926546812057
	pesos_i(867) := b"0000000000000000_0000000000000000_0001110010111111_1010011110100000"; -- 0.11229941993951797
	pesos_i(868) := b"1111111111111111_1111111111111111_1111010001001010_1110111001010000"; -- -0.045731645077466965
	pesos_i(869) := b"0000000000000000_0000000000000000_0010110111011001_0010011010000000"; -- 0.17909470200538635
	pesos_i(870) := b"1111111111111111_1111111111111111_1101101011000001_1001000101000000"; -- -0.14548389613628387
	pesos_i(871) := b"1111111111111111_1111111111111111_1010100110111100_1111101110000000"; -- -0.336960107088089
	pesos_i(872) := b"0000000000000000_0000000000000000_0010100100100011_0111010000000000"; -- 0.16069722175598145
	pesos_i(873) := b"0000000000000000_0000000000000000_0011001011110010_0101011001000000"; -- 0.19901026785373688
	pesos_i(874) := b"0000000000000000_0000000000000000_0000011100111111_0011111010001000"; -- 0.02830878086388111
	pesos_i(875) := b"0000000000000000_0000000000000000_0010101101100011_1001011100000000"; -- 0.16948837041854858
	pesos_i(876) := b"0000000000000000_0000000000000000_0010001110111011_0000001011000000"; -- 0.13957230746746063
	pesos_i(877) := b"0000000000000000_0000000000000000_0001111101010111_1010001000000000"; -- 0.12243092060089111
	pesos_i(878) := b"0000000000000000_0000000000000000_0001000101111011_1011110110100000"; -- 0.06829438358545303
	pesos_i(879) := b"1111111111111111_1111111111111111_1011011001011111_0010011110000000"; -- -0.28761056065559387
	pesos_i(880) := b"1111111111111111_1111111111111111_1001000011000100_0011101000000000"; -- -0.434505820274353
	pesos_i(881) := b"1111111111111111_1111111111111111_1000101100011000_0100110010000000"; -- -0.4566604793071747
	pesos_i(882) := b"0000000000000000_0000000000000000_0010010110011000_0000000011000000"; -- 0.14685063064098358
	pesos_i(883) := b"1111111111111111_1111111111111111_1010110111011001_0100011110000000"; -- -0.32090333104133606
	pesos_i(884) := b"1111111111111111_1111111111111111_1101110101011011_0000010001000000"; -- -0.1353299468755722
	pesos_i(885) := b"0000000000000000_0000000000000000_0011100011000111_0001010111000000"; -- 0.22178779542446136
	pesos_i(886) := b"1111111111111111_1111111111111111_1111111010001110_0110001011010110"; -- -0.00563986087217927
	pesos_i(887) := b"1111111111111111_1111111111111111_1011111100000001_0001001000000000"; -- -0.25388991832733154
	pesos_i(888) := b"1111111111111111_1111111111111111_1110000110001110_1101010011000000"; -- -0.11891432106494904
	pesos_i(889) := b"0000000000000000_0000000000000000_0101010101000000_1110100010000000"; -- 0.3330216705799103
	pesos_i(890) := b"1111111111111111_1111111111111111_1111111001011010_0101111011010010"; -- -0.006433557253330946
	pesos_i(891) := b"1111111111111111_1111111111111111_1111011110110110_1110001100000000"; -- -0.032365620136260986
	pesos_i(892) := b"0000000000000000_0000000000000000_0110011011011111_1110000100000000"; -- 0.40185362100601196
	pesos_i(893) := b"1111111111111111_1111111111111111_1110000101111101_1111110110100000"; -- -0.11917128413915634
	pesos_i(894) := b"1111111111111111_1111111111111111_1100011010010011_1000011110000000"; -- -0.22431138157844543
	pesos_i(895) := b"1111111111111111_1111111111111111_1011011101101101_1011011110000000"; -- -0.2834821045398712
	pesos_i(896) := b"0000000000000000_0000000000000000_0000011010100001_0010000111010000"; -- 0.025896180421113968
	pesos_i(897) := b"0000000000000000_0000000000000000_0001011101001101_1010110111000000"; -- 0.09102903306484222
	pesos_i(898) := b"1111111111111111_1111111111111111_1111100100111111_0000011110111000"; -- -0.02638198621571064
	pesos_i(899) := b"0000000000000000_0000000000000000_0010011101110101_1001110111000000"; -- 0.15413843095302582
	pesos_i(900) := b"1111111111111111_1111111111111111_1101100111001001_1000001001000000"; -- -0.1492689698934555
	pesos_i(901) := b"1111111111111111_1111111111111111_1100011101010110_1110110000000000"; -- -0.221329927444458
	pesos_i(902) := b"0000000000000000_0000000000000000_0011000101000010_0100110010000000"; -- 0.19241788983345032
	pesos_i(903) := b"0000000000000000_0000000000000000_0000110101010101_0111000111110000"; -- 0.052085038274526596
	pesos_i(904) := b"1111111111111111_1111111111111111_1011101101010010_0010101110000000"; -- -0.26827743649482727
	pesos_i(905) := b"1111111111111111_1111111111111111_1110010011011101_1010111100000000"; -- -0.1059923768043518
	pesos_i(906) := b"1111111111111111_1111111111111111_1100001010110001_1100100111000000"; -- -0.23947466909885406
	pesos_i(907) := b"1111111111111111_1111111111111111_1101100101111001_0001011100000000"; -- -0.15049606561660767
	pesos_i(908) := b"0000000000000000_0000000000000000_0000010001011111_0000101100100000"; -- 0.017075248062610626
	pesos_i(909) := b"0000000000000000_0000000000000000_0000011111101001_0111110001000000"; -- 0.030906453728675842
	pesos_i(910) := b"1111111111111111_1111111111111111_1110010101000110_0011011110100000"; -- -0.10439731925725937
	pesos_i(911) := b"1111111111111111_1111111111111111_1101101000011000_0001000000000000"; -- -0.1480703353881836
	pesos_i(912) := b"0000000000000000_0000000000000000_0000001100011011_1101110001011000"; -- 0.012143870815634727
	pesos_i(913) := b"0000000000000000_0000000000000000_0000110101110000_0010001011100000"; -- 0.05249231308698654
	pesos_i(914) := b"1111111111111111_1111111111111111_1110011000110001_1100010111000000"; -- -0.10080303251743317
	pesos_i(915) := b"1111111111111111_1111111111111111_1111111010011010_1111010011011100"; -- -0.005448051728308201
	pesos_i(916) := b"0000000000000000_0000000000000000_0001101110111100_1100111010100000"; -- 0.10834971815347672
	pesos_i(917) := b"1111111111111111_1111111111111111_1101100101111010_1000011010000000"; -- -0.1504741609096527
	pesos_i(918) := b"0000000000000000_0000000000000000_0000001111100101_0101000011000000"; -- 0.015217825770378113
	pesos_i(919) := b"1111111111111111_1111111111111111_1100110011000011_0111110011000000"; -- -0.20014210045337677
	pesos_i(920) := b"1111111111111111_1111111111111111_1001001111100010_0000111100000000"; -- -0.42233186960220337
	pesos_i(921) := b"1111111111111111_1111111111111111_1101100010010101_0101110101000000"; -- -0.1539708822965622
	pesos_i(922) := b"1111111111111111_1111111111111111_1110101000100001_0010010111000000"; -- -0.08543170988559723
	pesos_i(923) := b"0000000000000000_0000000000000000_0010010000000000_1111010101000000"; -- 0.14063961803913116
	pesos_i(924) := b"0000000000000000_0000000000000000_0010111000110100_0101100100000000"; -- 0.180486261844635
	pesos_i(925) := b"0000000000000000_0000000000000000_0011001100000010_0011011111000000"; -- 0.19925259053707123
	pesos_i(926) := b"0000000000000000_0000000000000000_0001110000011011_0111010110000000"; -- 0.10979399085044861
	pesos_i(927) := b"1111111111111111_1111111111111111_1110000000010011_0010001111100000"; -- -0.12470794469118118
	pesos_i(928) := b"0000000000000000_0000000000000000_0001100001001110_1011111101100000"; -- 0.09495159238576889
	pesos_i(929) := b"0000000000000000_0000000000000000_0000001101000101_1111011110000000"; -- 0.01278635859489441
	pesos_i(930) := b"0000000000000000_0000000000000000_0000010111001011_1111110100101000"; -- 0.02264387346804142
	pesos_i(931) := b"0000000000000000_0000000000000000_0000010100111101_0111010101000000"; -- 0.020469024777412415
	pesos_i(932) := b"0000000000000000_0000000000000000_0010000101011000_0001000110000000"; -- 0.13025006651878357
	pesos_i(933) := b"1111111111111111_1111111111111111_1111101000101000_0111101011111000"; -- -0.022819818928837776
	pesos_i(934) := b"1111111111111111_1111111111111111_1101000100010111_0000110010000000"; -- -0.1832420527935028
	pesos_i(935) := b"0000000000000000_0000000000000000_0010000110011100_0000110100000000"; -- 0.13128739595413208
	pesos_i(936) := b"0000000000000000_0000000000000000_0100010010011001_1000111100000000"; -- 0.2679681181907654
	pesos_i(937) := b"0000000000000000_0000000000000000_0100000101000011_1100100010000000"; -- 0.25494053959846497
	pesos_i(938) := b"1111111111111111_1111111111111111_1110110100011000_1101100101100000"; -- -0.07383958250284195
	pesos_i(939) := b"0000000000000000_0000000000000000_0001000101111000_1001000010100000"; -- 0.06824592500925064
	pesos_i(940) := b"1111111111111111_1111111111111111_1101000010010010_0100101001000000"; -- -0.18526779115200043
	pesos_i(941) := b"0000000000000000_0000000000000000_0000110111011000_0000011010010000"; -- 0.05407753959298134
	pesos_i(942) := b"1111111111111111_1111111111111111_1101111111100111_1011011011000000"; -- -0.1253705769777298
	pesos_i(943) := b"1111111111111111_1111111111111111_1111011111011010_1000011000000000"; -- -0.0318218469619751
	pesos_i(944) := b"1111111111111111_1111111111111111_1101100110011011_1101010010000000"; -- -0.14996597170829773
	pesos_i(945) := b"1111111111111111_1111111111111111_1110111101000111_0011110111000000"; -- -0.06531919538974762
	pesos_i(946) := b"1111111111111111_1111111111111111_1101010010000100_1101110100000000"; -- -0.16984766721725464
	pesos_i(947) := b"0000000000000000_0000000000000000_0000111011011100_1110011111110000"; -- 0.05805825814604759
	pesos_i(948) := b"1111111111111111_1111111111111111_1101101100010110_0010111000000000"; -- -0.14419281482696533
	pesos_i(949) := b"1111111111111111_1111111111111111_1011110100110100_0100011010000000"; -- -0.26092109084129333
	pesos_i(950) := b"0000000000000000_0000000000000000_0000110010010000_1100101100100000"; -- 0.04908437281847
	pesos_i(951) := b"1111111111111111_1111111111111111_1111010110111100_1001000010010000"; -- -0.04009148105978966
	pesos_i(952) := b"1111111111111111_1111111111111111_1100001101011000_1110110101000000"; -- -0.23692433536052704
	pesos_i(953) := b"0000000000000000_0000000000000000_0100000111100011_0100111100000000"; -- 0.25737470388412476
	pesos_i(954) := b"1111111111111111_1111111111111111_1101100010101010_0000101100000000"; -- -0.15365535020828247
	pesos_i(955) := b"0000000000000000_0000000000000000_0011011011100010_0110000111000000"; -- 0.2143918126821518
	pesos_i(956) := b"0000000000000000_0000000000000000_0000101101000100_1010000101000000"; -- 0.04401595890522003
	pesos_i(957) := b"0000000000000000_0000000000000000_0001110111100010_1011100001100000"; -- 0.11674072593450546
	pesos_i(958) := b"0000000000000000_0000000000000000_0011101101000000_0010010001000000"; -- 0.2314474731683731
	pesos_i(959) := b"0000000000000000_0000000000000000_0000011110100000_1010110110111000"; -- 0.029795510694384575
	pesos_i(960) := b"0000000000000000_0000000000000000_0011001011011110_0111110111000000"; -- 0.1987074464559555
	pesos_i(961) := b"1111111111111111_1111111111111111_1100101110001001_0101011011000000"; -- -0.20493562519550323
	pesos_i(962) := b"1111111111111111_1111111111111111_1110101011010001_1001001111000000"; -- -0.08273960649967194
	pesos_i(963) := b"0000000000000000_0000000000000000_0000001100110110_0111101001001000"; -- 0.01255001313984394
	pesos_i(964) := b"1111111111111111_1111111111111111_1010111000101111_1011000010000000"; -- -0.31958481669425964
	pesos_i(965) := b"0000000000000000_0000000000000000_0010010011101100_0011101101000000"; -- 0.14422960579395294
	pesos_i(966) := b"0000000000000000_0000000000000000_0001110101101101_0100001010100000"; -- 0.11494842916727066
	pesos_i(967) := b"1111111111111111_1111111111111111_1100000110100110_1001010000000000"; -- -0.24355196952819824
	pesos_i(968) := b"0000000000000000_0000000000000000_0001100010110100_0011010010000000"; -- 0.09649971127510071
	pesos_i(969) := b"1111111111111111_1111111111111111_1101011000010000_1011000010000000"; -- -0.16380783915519714
	pesos_i(970) := b"0000000000000000_0000000000000000_0100111000110010_0100111100000000"; -- 0.30545514822006226
	pesos_i(971) := b"0000000000000000_0000000000000000_0000100011110110_1111110111010000"; -- 0.035018790513277054
	pesos_i(972) := b"0000000000000000_0000000000000000_0000001100000100_0000110001000000"; -- 0.011780515313148499
	pesos_i(973) := b"0000000000000000_0000000000000000_0001010011111111_0001000001000000"; -- 0.0820169597864151
	pesos_i(974) := b"1111111111111111_1111111111111111_1110011101111000_0000010010100000"; -- -0.09582491964101791
	pesos_i(975) := b"1111111111111111_1111111111111111_1110011111101010_1100101100100000"; -- -0.094073586165905
	pesos_i(976) := b"1111111111111111_1111111111111111_1101000001010100_0101100111000000"; -- -0.1862129122018814
	pesos_i(977) := b"0000000000000000_0000000000000000_0000101110010110_0101101011110000"; -- 0.04526298865675926
	pesos_i(978) := b"1111111111111111_1111111111111111_1111100110111001_0011111001010000"; -- -0.024517159909009933
	pesos_i(979) := b"0000000000000000_0000000000000000_0001110011010011_1011110011000000"; -- 0.11260585486888885
	pesos_i(980) := b"1111111111111111_1111111111111111_1111111110111001_1001100110101001"; -- -0.0010742151644080877
	pesos_i(981) := b"1111111111111111_1111111111111111_1011111110000111_0101111000000000"; -- -0.2518407106399536
	pesos_i(982) := b"1111111111111111_1111111111111111_1100011111000001_1000110011000000"; -- -0.21970291435718536
	pesos_i(983) := b"1111111111111111_1111111111111111_1110001110111100_1111111011000000"; -- -0.11039741337299347
	pesos_i(984) := b"0000000000000000_0000000000000000_0001010100110110_1100111011100000"; -- 0.08286755532026291
	pesos_i(985) := b"0000000000000000_0000000000000000_0011011011000101_1010001101000000"; -- 0.21395321190357208
	pesos_i(986) := b"1111111111111111_1111111111111111_1110010001101111_1110001111000000"; -- -0.1076676994562149
	pesos_i(987) := b"1111111111111111_1111111111111111_1011011110100111_0011111100000000"; -- -0.28260427713394165
	pesos_i(988) := b"0000000000000000_0000000000000000_0011110010011000_1010000001000000"; -- 0.23670388758182526
	pesos_i(989) := b"1111111111111111_1111111111111111_1100100011010100_0111110001000000"; -- -0.21550773084163666
	pesos_i(990) := b"0000000000000000_0000000000000000_0000011111000111_1001100110110000"; -- 0.030389409512281418
	pesos_i(991) := b"0000000000000000_0000000000000000_0000101001001111_0101001110100000"; -- 0.04027292877435684
	pesos_i(992) := b"1111111111111111_1111111111111111_1111001101101110_0000100110110000"; -- -0.04910220578312874
	pesos_i(993) := b"1111111111111111_1111111111111111_1111001111010100_0010111100000000"; -- -0.04754358530044556
	pesos_i(994) := b"1111111111111111_1111111111111111_1110110100001010_1101101100000000"; -- -0.07405310869216919
	pesos_i(995) := b"1111111111111111_1111111111111111_1111111110010101_0101010000010101"; -- -0.0016276787500828505
	pesos_i(996) := b"0000000000000000_0000000000000000_0010010110000000_1001001111000000"; -- 0.14649318158626556
	pesos_i(997) := b"0000000000000000_0000000000000000_0000100100011000_1100100000000000"; -- 0.03553438186645508
	pesos_i(998) := b"0000000000000000_0000000000000000_0001010010010000_1000000010100000"; -- 0.08032993227243423
	pesos_i(999) := b"1111111111111111_1111111111111111_1010111100101010_1110000100000000"; -- -0.31575196981430054
	pesos_i(1000) := b"1111111111111111_1111111111111111_1101101100001001_1101010011000000"; -- -0.14438124001026154
	pesos_i(1001) := b"0000000000000000_0000000000000000_0010011111111101_1001110001000000"; -- 0.15621353685855865
	pesos_i(1002) := b"0000000000000000_0000000000000000_0010010011011001_0110000111000000"; -- 0.1439419835805893
	pesos_i(1003) := b"0000000000000000_0000000000000000_0100011101100101_1011001100000000"; -- 0.2788955569267273
	pesos_i(1004) := b"1111111111111111_1111111111111111_1111101000111111_0000011111100000"; -- -0.022475726902484894
	pesos_i(1005) := b"1111111111111111_1111111111111111_1111011110011000_1001111001100000"; -- -0.0328274741768837
	pesos_i(1006) := b"0000000000000000_0000000000000000_0010110010110100_0110101111000000"; -- 0.17462800443172455
	pesos_i(1007) := b"1111111111111111_1111111111111111_1110010110111111_0110000000100000"; -- -0.10254859179258347
	pesos_i(1008) := b"1111111111111111_1111111111111111_1110000110010000_1011100101000000"; -- -0.11888544261455536
	pesos_i(1009) := b"1111111111111111_1111111111111111_1100101111101010_0001000001000000"; -- -0.2034597247838974
	pesos_i(1010) := b"0000000000000000_0000000000000000_0001000110111000_0010010111100000"; -- 0.06921612471342087
	pesos_i(1011) := b"1111111111111111_1111111111111111_1100101110101000_1010011101000000"; -- -0.20445780456066132
	pesos_i(1012) := b"1111111111111111_1111111111111111_1101101110110011_0110111100000000"; -- -0.14179331064224243
	pesos_i(1013) := b"0000000000000000_0000000000000000_0010011111010001_0011101100000000"; -- 0.15553635358810425
	pesos_i(1014) := b"0000000000000000_0000000000000000_0001100110001111_1111010001100000"; -- 0.09985282272100449
	pesos_i(1015) := b"1111111111111111_1111111111111111_1100001011110100_0111011011000000"; -- -0.23845727741718292
	pesos_i(1016) := b"0000000000000000_0000000000000000_0000100111100000_0100001110010000"; -- 0.03857824578881264
	pesos_i(1017) := b"0000000000000000_0000000000000000_0000100100110000_0011001100010000"; -- 0.03589171543717384
	pesos_i(1018) := b"0000000000000000_0000000000000000_0011000010001001_0001111000000000"; -- 0.18959224224090576
	pesos_i(1019) := b"1111111111111111_1111111111111111_1011110011001010_0110000100000000"; -- -0.2625369429588318
	pesos_i(1020) := b"1111111111111111_1111111111111111_1111001010001010_0100000111100000"; -- -0.05257786065340042
	pesos_i(1021) := b"1111111111111111_1111111111111111_1111111010011110_0110110100010010"; -- -0.005395110230892897
	pesos_i(1022) := b"1111111111111111_1111111111111111_1101110101011000_0110001000000000"; -- -0.135370135307312
	pesos_i(1023) := b"0000000000000000_0000000000000000_0001000100010100_1111100000000000"; -- 0.0667262077331543
	pesos_i(1024) := b"1111111111111111_1111111111111111_1110110100110001_1010010000100000"; -- -0.07346128672361374
	pesos_i(1025) := b"1111111111111111_1111111111111111_1110101011100001_0111000010000000"; -- -0.08249756693840027
	pesos_i(1026) := b"1111111111111111_1111111111111111_1111100011010010_0001010000011000"; -- -0.028044456616044044
	pesos_i(1027) := b"1111111111111111_1111111111111111_1111111110000110_1101010101101001"; -- -0.0018488520290702581
	pesos_i(1028) := b"1111111111111111_1111111111111111_1111000001110010_0001111111110000"; -- -0.060758594423532486
	pesos_i(1029) := b"1111111111111111_1111111111111111_1110110001101010_0110110010100000"; -- -0.07650109380483627
	pesos_i(1030) := b"0000000000000000_0000000000000000_0011101110100001_1100010000000000"; -- 0.23293709754943848
	pesos_i(1031) := b"0000000000000000_0000000000000000_0011010111010110_0111001000000000"; -- 0.2103034257888794
	pesos_i(1032) := b"0000000000000000_0000000000000000_0010110111001001_0011000101000000"; -- 0.1788512021303177
	pesos_i(1033) := b"1111111111111111_1111111111111111_1111100111100111_0001001101001000"; -- -0.023817820474505424
	pesos_i(1034) := b"0000000000000000_0000000000000000_0000101110100010_0010011101100000"; -- 0.04544302076101303
	pesos_i(1035) := b"0000000000000000_0000000000000000_0010001010101111_0001110000000000"; -- 0.1354844570159912
	pesos_i(1036) := b"0000000000000000_0000000000000000_0001010001000111_1000100011000000"; -- 0.07921652495861053
	pesos_i(1037) := b"1111111111111111_1111111111111111_1111001010100110_0101110110010000"; -- -0.0521489642560482
	pesos_i(1038) := b"0000000000000000_0000000000000000_0011010110100001_0000001110000000"; -- 0.2094881236553192
	pesos_i(1039) := b"0000000000000000_0000000000000000_0001100011001110_1001010111100000"; -- 0.09690224379301071
	pesos_i(1040) := b"1111111111111111_1111111111111111_1111111000000101_1110111101011100"; -- -0.0077219391241669655
	pesos_i(1041) := b"0000000000000000_0000000000000000_0000011000001101_0000110011010000"; -- 0.023636627942323685
	pesos_i(1042) := b"0000000000000000_0000000000000000_0010100110110101_0101001100000000"; -- 0.16292303800582886
	pesos_i(1043) := b"0000000000000000_0000000000000000_0001100110100110_1010101111000000"; -- 0.10019944608211517
	pesos_i(1044) := b"1111111111111111_1111111111111111_1100100101110001_0000111011000000"; -- -0.21311862766742706
	pesos_i(1045) := b"0000000000000000_0000000000000000_0010010011111011_0001101101000000"; -- 0.14445658028125763
	pesos_i(1046) := b"0000000000000000_0000000000000000_0001001010010001_0100010010100000"; -- 0.07252911478281021
	pesos_i(1047) := b"1111111111111111_1111111111111111_1100001110100100_1001001100000000"; -- -0.23577004671096802
	pesos_i(1048) := b"1111111111111111_1111111111111111_1101001010100101_1001111001000000"; -- -0.1771603673696518
	pesos_i(1049) := b"1111111111111111_1111111111111111_1110000110010001_0001110110100000"; -- -0.11887945979833603
	pesos_i(1050) := b"0000000000000000_0000000000000000_0011011010011100_0011100110000000"; -- 0.21332129836082458
	pesos_i(1051) := b"0000000000000000_0000000000000000_0000101010110001_0110000011000000"; -- 0.04176907241344452
	pesos_i(1052) := b"0000000000000000_0000000000000000_0001111100111011_1011101101100000"; -- 0.12200518697500229
	pesos_i(1053) := b"1111111111111111_1111111111111111_1100100000100000_0000111111000000"; -- -0.2182607799768448
	pesos_i(1054) := b"0000000000000000_0000000000000000_0001100110110011_1010001011100000"; -- 0.10039728134870529
	pesos_i(1055) := b"1111111111111111_1111111111111111_1100100000100110_1101001001000000"; -- -0.21815763413906097
	pesos_i(1056) := b"1111111111111111_1111111111111111_1100101101110000_1011001111000000"; -- -0.20531155169010162
	pesos_i(1057) := b"0000000000000000_0000000000000000_0000111001001100_0111100011010000"; -- 0.05585436895489693
	pesos_i(1058) := b"0000000000000000_0000000000000000_0000011001000010_0011101100110000"; -- 0.024448107928037643
	pesos_i(1059) := b"1111111111111111_1111111111111111_1111010111100011_1101100111000000"; -- -0.03949202597141266
	pesos_i(1060) := b"0000000000000000_0000000000000000_0001001110101111_1000101001000000"; -- 0.0768972784280777
	pesos_i(1061) := b"0000000000000000_0000000000000000_0010011110110101_0001100110000000"; -- 0.15510711073875427
	pesos_i(1062) := b"1111111111111111_1111111111111111_1100011001011100_1000101001000000"; -- -0.2251504510641098
	pesos_i(1063) := b"0000000000000000_0000000000000000_0001110011111001_1110011111100000"; -- 0.1131882593035698
	pesos_i(1064) := b"0000000000000000_0000000000000000_0011000001100011_1001010100000000"; -- 0.18901950120925903
	pesos_i(1065) := b"0000000000000000_0000000000000000_0010100000001001_1000010101000000"; -- 0.15639527142047882
	pesos_i(1066) := b"0000000000000000_0000000000000000_0010010001100000_1010111000000000"; -- 0.14210021495819092
	pesos_i(1067) := b"1111111111111111_1111111111111111_1110101000000101_1010110111100000"; -- -0.08585084229707718
	pesos_i(1068) := b"0000000000000000_0000000000000000_0010011101100111_1100000100000000"; -- 0.15392690896987915
	pesos_i(1069) := b"0000000000000000_0000000000000000_0010100011011111_0101000011000000"; -- 0.1596575230360031
	pesos_i(1070) := b"0000000000000000_0000000000000000_0000011100001000_1010111100011000"; -- 0.02747625671327114
	pesos_i(1071) := b"0000000000000000_0000000000000000_0010110101010011_1000101111000000"; -- 0.17705605924129486
	pesos_i(1072) := b"0000000000000000_0000000000000000_0010111110000010_1101001110000000"; -- 0.185589998960495
	pesos_i(1073) := b"1111111111111111_1111111111111111_1110011101001010_0000001010100000"; -- -0.09652694314718246
	pesos_i(1074) := b"1111111111111111_1111111111111111_1111011101010111_1101101110110000"; -- -0.033815640956163406
	pesos_i(1075) := b"1111111111111111_1111111111111111_1111010111110111_0111010000000000"; -- -0.039192914962768555
	pesos_i(1076) := b"1111111111111111_1111111111111111_1101011100011010_0110011100000000"; -- -0.15975338220596313
	pesos_i(1077) := b"0000000000000000_0000000000000000_0000000110001111_0100110001101010"; -- 0.006092811468988657
	pesos_i(1078) := b"1111111111111111_1111111111111111_1101001001100000_1100000100000000"; -- -0.17821115255355835
	pesos_i(1079) := b"0000000000000000_0000000000000000_0011001110011001_1001100010000000"; -- 0.20156243443489075
	pesos_i(1080) := b"1111111111111111_1111111111111111_1111100110110110_1000010111000000"; -- -0.02455867826938629
	pesos_i(1081) := b"0000000000000000_0000000000000000_0000101011101000_1111000010100000"; -- 0.04261688143014908
	pesos_i(1082) := b"1111111111111111_1111111111111111_1100100011101100_0111001001000000"; -- -0.2151421159505844
	pesos_i(1083) := b"0000000000000000_0000000000000000_0000001110101011_0011000110011100"; -- 0.014330959878861904
	pesos_i(1084) := b"0000000000000000_0000000000000000_0010101000111011_1110000110000000"; -- 0.16497620940208435
	pesos_i(1085) := b"1111111111111111_1111111111111111_1100100000100100_0010010101000000"; -- -0.21819846332073212
	pesos_i(1086) := b"0000000000000000_0000000000000000_0001111001110110_0001011000000000"; -- 0.11898934841156006
	pesos_i(1087) := b"0000000000000000_0000000000000000_0000001000001011_0000011011001100"; -- 0.007980751805007458
	pesos_i(1088) := b"0000000000000000_0000000000000000_0010100010111001_1000101000000000"; -- 0.1590811014175415
	pesos_i(1089) := b"0000000000000000_0000000000000000_0001111110001010_1010110011100000"; -- 0.12320976704359055
	pesos_i(1090) := b"1111111111111111_1111111111111111_1111110011110000_0011100100001000"; -- -0.011959491297602654
	pesos_i(1091) := b"0000000000000000_0000000000000000_0010000000011111_1011101000000000"; -- 0.12548410892486572
	pesos_i(1092) := b"0000000000000000_0000000000000000_0001010011100101_1011101000100000"; -- 0.08163035660982132
	pesos_i(1093) := b"0000000000000000_0000000000000000_0000111111001011_0101111110100000"; -- 0.06169698387384415
	pesos_i(1094) := b"0000000000000000_0000000000000000_0000011001001011_1000011111111000"; -- 0.024590013548731804
	pesos_i(1095) := b"1111111111111111_1111111111111111_1111101010000100_1011111110010000"; -- -0.021411921828985214
	pesos_i(1096) := b"1111111111111111_1111111111111111_1111001111101010_1000000100010000"; -- -0.047203000634908676
	pesos_i(1097) := b"0000000000000000_0000000000000000_0000011100100101_1101011010100000"; -- 0.027921117842197418
	pesos_i(1098) := b"1111111111111111_1111111111111111_1111011011011100_1011111011000000"; -- -0.035694196820259094
	pesos_i(1099) := b"0000000000000000_0000000000000000_0000110110111110_0110110100100000"; -- 0.053686924278736115
	pesos_i(1100) := b"0000000000000000_0000000000000000_0010001111101111_0110111010000000"; -- 0.14037218689918518
	pesos_i(1101) := b"0000000000000000_0000000000000000_0000011100010000_0100110111011000"; -- 0.027592530474066734
	pesos_i(1102) := b"1111111111111111_1111111111111111_1011100010110100_0001010010000000"; -- -0.2785021960735321
	pesos_i(1103) := b"0000000000000000_0000000000000000_0010110100001001_0001000011000000"; -- 0.1759195774793625
	pesos_i(1104) := b"1111111111111111_1111111111111111_1111011110111011_0001110101110000"; -- -0.032301101833581924
	pesos_i(1105) := b"0000000000000000_0000000000000000_0000001010100110_1111001101101100"; -- 0.010359968058764935
	pesos_i(1106) := b"1111111111111111_1111111111111111_1111101011111111_1001000100100000"; -- -0.01953785866498947
	pesos_i(1107) := b"1111111111111111_1111111111111111_1101001010011111_0101000010000000"; -- -0.17725655436515808
	pesos_i(1108) := b"1111111111111111_1111111111111111_1101100001100101_1001001011000000"; -- -0.1547001153230667
	pesos_i(1109) := b"0000000000000000_0000000000000000_0000100011111101_1000101111110000"; -- 0.035118814557790756
	pesos_i(1110) := b"1111111111111111_1111111111111111_1111000110101011_1111001010010000"; -- -0.05597003921866417
	pesos_i(1111) := b"0000000000000000_0000000000000000_0010111010111100_0101010111000000"; -- 0.1825612634420395
	pesos_i(1112) := b"0000000000000000_0000000000000000_0011011011010010_1000010111000000"; -- 0.2141498178243637
	pesos_i(1113) := b"1111111111111111_1111111111111111_1111100100000010_1101011101010000"; -- -0.0273003987967968
	pesos_i(1114) := b"1111111111111111_1111111111111111_1100000111101111_0100101000000000"; -- -0.24244248867034912
	pesos_i(1115) := b"0000000000000000_0000000000000000_0001111000000001_1101110110100000"; -- 0.11721596866846085
	pesos_i(1116) := b"0000000000000000_0000000000000000_0001001111001001_0100011111100000"; -- 0.07729005068540573
	pesos_i(1117) := b"1111111111111111_1111111111111111_1111010000111101_1100110100010000"; -- -0.045931991189718246
	pesos_i(1118) := b"0000000000000000_0000000000000000_0000001111110011_1010110010011000"; -- 0.015436923131346703
	pesos_i(1119) := b"1111111111111111_1111111111111111_1110100001110001_0110010110000000"; -- -0.0920197069644928
	pesos_i(1120) := b"1111111111111111_1111111111111111_1101110101110010_1010101011000000"; -- -0.1349690705537796
	pesos_i(1121) := b"1111111111111111_1111111111111111_1111101001111011_1011101010000000"; -- -0.02154955267906189
	pesos_i(1122) := b"1111111111111111_1111111111111111_1110110000011000_1101010011000000"; -- -0.07774610817432404
	pesos_i(1123) := b"1111111111111111_1111111111111111_1110110101000101_1110011111000000"; -- -0.0731520801782608
	pesos_i(1124) := b"1111111111111111_1111111111111111_1101011101111001_1011010011000000"; -- -0.15829916298389435
	pesos_i(1125) := b"0000000000000000_0000000000000000_0001101001111100_0110100011000000"; -- 0.10346083343029022
	pesos_i(1126) := b"0000000000000000_0000000000000000_0010011000001011_1101111111000000"; -- 0.148618683218956
	pesos_i(1127) := b"0000000000000000_0000000000000000_0000101011010000_0100100111010000"; -- 0.042240727692842484
	pesos_i(1128) := b"1111111111111111_1111111111111111_1001111100101110_0000010100000000"; -- -0.3782040476799011
	pesos_i(1129) := b"0000000000000000_0000000000000000_0010010100001011_0001010001000000"; -- 0.1447003036737442
	pesos_i(1130) := b"1111111111111111_1111111111111111_1011101000011001_0010001110000000"; -- -0.273053914308548
	pesos_i(1131) := b"1111111111111111_1111111111111111_1111000001011100_1111000000110000"; -- -0.06108187511563301
	pesos_i(1132) := b"0000000000000000_0000000000000000_0000000000111100_0101110011100100"; -- 0.0009210639400407672
	pesos_i(1133) := b"1111111111111111_1111111111111111_1101110110000111_1101000110000000"; -- -0.13464632630348206
	pesos_i(1134) := b"0000000000000000_0000000000000000_0001011111000000_0101110000000000"; -- 0.09277892112731934
	pesos_i(1135) := b"1111111111111111_1111111111111111_1110011101101111_0010000001100000"; -- -0.0959605947136879
	pesos_i(1136) := b"1111111111111111_1111111111111111_1110010110011010_0001010101100000"; -- -0.10311762243509293
	pesos_i(1137) := b"1111111111111111_1111111111111111_1010111010000100_0010110000000000"; -- -0.3182957172393799
	pesos_i(1138) := b"1111111111111111_1111111111111111_1111100100001111_1100110011011000"; -- -0.02710265852510929
	pesos_i(1139) := b"1111111111111111_1111111111111111_1111010001100000_0111100001110000"; -- -0.045402977615594864
	pesos_i(1140) := b"1111111111111111_1111111111111111_1100001111001110_0001001101000000"; -- -0.23513679206371307
	pesos_i(1141) := b"0000000000000000_0000000000000000_0000010101111010_1100000000001000"; -- 0.021404268220067024
	pesos_i(1142) := b"1111111111111111_1111111111111111_1111011111010011_1001001110100000"; -- -0.03192784637212753
	pesos_i(1143) := b"0000000000000000_0000000000000000_0011100111111010_0000001010000000"; -- 0.22647109627723694
	pesos_i(1144) := b"1111111111111111_1111111111111111_1111100001001001_0001110110011000"; -- -0.03013434447348118
	pesos_i(1145) := b"0000000000000000_0000000000000000_0011011111111001_1010100100000000"; -- 0.21865326166152954
	pesos_i(1146) := b"0000000000000000_0000000000000000_0000001100111100_0001000011010100"; -- 0.012635280378162861
	pesos_i(1147) := b"0000000000000000_0000000000000000_0000110101001001_0011001001100000"; -- 0.05189814418554306
	pesos_i(1148) := b"1111111111111111_1111111111111111_1100101110000100_0100100101000000"; -- -0.2050127238035202
	pesos_i(1149) := b"1111111111111111_1111111111111111_1111110100101110_0111001010001000"; -- -0.011010019108653069
	pesos_i(1150) := b"1111111111111111_1111111111111111_1101110110100010_1101010100000000"; -- -0.13423413038253784
	pesos_i(1151) := b"1111111111111111_1111111111111111_1110011110100010_1010111000000000"; -- -0.09517395496368408
	pesos_i(1152) := b"0000000000000000_0000000000000000_0011101111110110_0000111100000000"; -- 0.23422330617904663
	pesos_i(1153) := b"0000000000000000_0000000000000000_0001111100110110_1011010011100000"; -- 0.12192850559949875
	pesos_i(1154) := b"0000000000000000_0000000000000000_0010001111000000_0011101111000000"; -- 0.13965199887752533
	pesos_i(1155) := b"1111111111111111_1111111111111111_1101101001110100_1101010110000000"; -- -0.14665475487709045
	pesos_i(1156) := b"1111111111111111_1111111111111111_1101101111010100_0001111001000000"; -- -0.14129458367824554
	pesos_i(1157) := b"1111111111111111_1111111111111111_1010111011010001_0110111110000000"; -- -0.31711676716804504
	pesos_i(1158) := b"0000000000000000_0000000000000000_0000001011111110_0110010000110100"; -- 0.011694204993546009
	pesos_i(1159) := b"0000000000000000_0000000000000000_0010001111010010_1101101100000000"; -- 0.1399361491203308
	pesos_i(1160) := b"0000000000000000_0000000000000000_0001000110011000_1000001010100000"; -- 0.06873337179422379
	pesos_i(1161) := b"1111111111111111_1111111111111111_1100000111101110_1000111111000000"; -- -0.24245359003543854
	pesos_i(1162) := b"1111111111111111_1111111111111111_1110101011000101_0001110010100000"; -- -0.0829298123717308
	pesos_i(1163) := b"0000000000000000_0000000000000000_0001010000011100_1101100001000000"; -- 0.07856513559818268
	pesos_i(1164) := b"0000000000000000_0000000000000000_0000000100111011_1010111111100100"; -- 0.0048170024529099464
	pesos_i(1165) := b"1111111111111111_1111111111111111_1110100110110010_1010111010100000"; -- -0.0871172770857811
	pesos_i(1166) := b"0000000000000000_0000000000000000_0011000001001111_0110001100000000"; -- 0.18871134519577026
	pesos_i(1167) := b"0000000000000000_0000000000000000_0010001001100010_1010001111000000"; -- 0.13431762158870697
	pesos_i(1168) := b"1111111111111111_1111111111111111_1011111010001010_1110111000000000"; -- -0.25569260120391846
	pesos_i(1169) := b"1111111111111111_1111111111111111_1111101010110111_1000101100100000"; -- -0.020636849105358124
	pesos_i(1170) := b"1111111111111111_1111111111111111_1001110101000111_0011011000000000"; -- -0.38563215732574463
	pesos_i(1171) := b"0000000000000000_0000000000000000_0000000010101110_1111110001110000"; -- 0.0026700757443904877
	pesos_i(1172) := b"1111111111111111_1111111111111111_1111011001001110_0110110101100000"; -- -0.03786579519510269
	pesos_i(1173) := b"0000000000000000_0000000000000000_0010010010111101_1010000011000000"; -- 0.14351849257946014
	pesos_i(1174) := b"0000000000000000_0000000000000000_0001111111111111_1011000101100000"; -- 0.12499531358480453
	pesos_i(1175) := b"0000000000000000_0000000000000000_0001000101100101_1000011101000000"; -- 0.06795544922351837
	pesos_i(1176) := b"1111111111111111_1111111111111111_1100000011110110_1000010101000000"; -- -0.24623839557170868
	pesos_i(1177) := b"0000000000000000_0000000000000000_0001111010010001_0001010010000000"; -- 0.1194012463092804
	pesos_i(1178) := b"0000000000000000_0000000000000000_0001000011111011_0011110101000000"; -- 0.06633360683917999
	pesos_i(1179) := b"1111111111111111_1111111111111111_1111001111000011_1101000010010000"; -- -0.04779335483908653
	pesos_i(1180) := b"1111111111111111_1111111111111111_1100011110110011_1010011100000000"; -- -0.219914972782135
	pesos_i(1181) := b"1111111111111111_1111111111111111_1110011100101001_1010011100000000"; -- -0.09702068567276001
	pesos_i(1182) := b"0000000000000000_0000000000000000_0001101100001110_1011010100000000"; -- 0.10569316148757935
	pesos_i(1183) := b"0000000000000000_0000000000000000_0000000011110010_1110001101100001"; -- 0.003706179792061448
	pesos_i(1184) := b"1111111111111111_1111111111111111_1101001011111000_0000110011000000"; -- -0.1759025603532791
	pesos_i(1185) := b"1111111111111111_1111111111111111_1111001000100100_1100110001000000"; -- -0.054126009345054626
	pesos_i(1186) := b"0000000000000000_0000000000000000_0011110010110001_0101111010000000"; -- 0.23708143830299377
	pesos_i(1187) := b"1111111111111111_1111111111111111_1110111011010000_0100100000100000"; -- -0.06713437288999557
	pesos_i(1188) := b"1111111111111111_1111111111111111_1101100101001001_0100010100000000"; -- -0.151225745677948
	pesos_i(1189) := b"1111111111111111_1111111111111111_1111101010011010_1000001111011000"; -- -0.021079787984490395
	pesos_i(1190) := b"1111111111111111_1111111111111111_1111110000001100_0111010110110000"; -- -0.015434879809617996
	pesos_i(1191) := b"1111111111111111_1111111111111111_1101100001010010_0010000101000000"; -- -0.15499679744243622
	pesos_i(1192) := b"1111111111111111_1111111111111111_1111000000001101_1011100001110000"; -- -0.06229064241051674
	pesos_i(1193) := b"1111111111111111_1111111111111111_1100101000100010_1011011110000000"; -- -0.21040776371955872
	pesos_i(1194) := b"0000000000000000_0000000000000000_0010001000010111_1011100010000000"; -- 0.13317444920539856
	pesos_i(1195) := b"1111111111111111_1111111111111111_1110110001000011_1011101001000000"; -- -0.07709155976772308
	pesos_i(1196) := b"1111111111111111_1111111111111111_1111010110000100_0101111101100000"; -- -0.04094890505075455
	pesos_i(1197) := b"1111111111111111_1111111111111111_1110100100110101_1100101001100000"; -- -0.08902297168970108
	pesos_i(1198) := b"0000000000000000_0000000000000000_0000011100101101_1001001100100000"; -- 0.02803916484117508
	pesos_i(1199) := b"1111111111111111_1111111111111111_1101101011000111_1111010100000000"; -- -0.14538639783859253
	pesos_i(1200) := b"1111111111111111_1111111111111111_1110110000100111_0000101100100000"; -- -0.07752924412488937
	pesos_i(1201) := b"0000000000000000_0000000000000000_0010110101010000_1110111000000000"; -- 0.17701613903045654
	pesos_i(1202) := b"0000000000000000_0000000000000000_0000100011010101_0101100111000000"; -- 0.03450547158718109
	pesos_i(1203) := b"1111111111111111_1111111111111111_1110101111000010_1010101000000000"; -- -0.07906091213226318
	pesos_i(1204) := b"0000000000000000_0000000000000000_0001100101100000_0011100010100000"; -- 0.0991244688630104
	pesos_i(1205) := b"1111111111111111_1111111111111111_1111011111001000_1010001000010000"; -- -0.03209483250975609
	pesos_i(1206) := b"0000000000000000_0000000000000000_0000001000011010_1110101111011000"; -- 0.008223285898566246
	pesos_i(1207) := b"0000000000000000_0000000000000000_0011011101111000_1011110100000000"; -- 0.21668606996536255
	pesos_i(1208) := b"0000000000000000_0000000000000000_0000001001000100_1000000110010000"; -- 0.008857820183038712
	pesos_i(1209) := b"0000000000000000_0000000000000000_0000011001011111_0100100111111000"; -- 0.02489149384200573
	pesos_i(1210) := b"1111111111111111_1111111111111111_1111000111001000_1011011011000000"; -- -0.0555310994386673
	pesos_i(1211) := b"0000000000000000_0000000000000000_0010101000100011_1101101111000000"; -- 0.1646096557378769
	pesos_i(1212) := b"0000000000000000_0000000000000000_0010000001011111_1111100011000000"; -- 0.12646441161632538
	pesos_i(1213) := b"1111111111111111_1111111111111111_1001100001000011_0010000010000000"; -- -0.4052257239818573
	pesos_i(1214) := b"0000000000000000_0000000000000000_0001111011101101_0101010011100000"; -- 0.12080889195203781
	pesos_i(1215) := b"1111111111111111_1111111111111111_1111100001010100_0100000001111000"; -- -0.029964419081807137
	pesos_i(1216) := b"1111111111111111_1111111111111111_1100110001101010_1101001011000000"; -- -0.2014950066804886
	pesos_i(1217) := b"1111111111111111_1111111111111111_1110111001111111_1010110010100000"; -- -0.06836434453725815
	pesos_i(1218) := b"0000000000000000_0000000000000000_0000110111001010_0100101011010000"; -- 0.05386798456311226
	pesos_i(1219) := b"0000000000000000_0000000000000000_0001000110011111_1011111010000000"; -- 0.06884375214576721
	pesos_i(1220) := b"0000000000000000_0000000000000000_0010100111111011_0100000010000000"; -- 0.1639900505542755
	pesos_i(1221) := b"0000000000000000_0000000000000000_0001010011001011_0101001010000000"; -- 0.08122745156288147
	pesos_i(1222) := b"0000000000000000_0000000000000000_0101100001011000_1010111110000000"; -- 0.3451032340526581
	pesos_i(1223) := b"0000000000000000_0000000000000000_0000011100001101_1111100100001000"; -- 0.02755695767700672
	pesos_i(1224) := b"0000000000000000_0000000000000000_0010110011010001_0010010110000000"; -- 0.17506632208824158
	pesos_i(1225) := b"1111111111111111_1111111111111111_1110100100000000_0111100010100000"; -- -0.08983656018972397
	pesos_i(1226) := b"0000000000000000_0000000000000000_0011001110100110_1100001110000000"; -- 0.2017633616924286
	pesos_i(1227) := b"0000000000000000_0000000000000000_0100010011011101_0000100100000000"; -- 0.2689977288246155
	pesos_i(1228) := b"1111111111111111_1111111111111111_1011010110101101_1011001010000000"; -- -0.2903183400630951
	pesos_i(1229) := b"1111111111111111_1111111111111111_1111010110011000_0111101100000000"; -- -0.04064208269119263
	pesos_i(1230) := b"1111111111111111_1111111111111111_1011010011100001_0100110000000000"; -- -0.29343724250793457
	pesos_i(1231) := b"1111111111111111_1111111111111111_1111101010010011_1010100000100000"; -- -0.021184436976909637
	pesos_i(1232) := b"0000000000000000_0000000000000000_0001010110010001_1001100010000000"; -- 0.08425286412239075
	pesos_i(1233) := b"0000000000000000_0000000000000000_0001000010101011_1011101001100000"; -- 0.06512036174535751
	pesos_i(1234) := b"0000000000000000_0000000000000000_0000100110100100_1110001000010000"; -- 0.03767216578125954
	pesos_i(1235) := b"1111111111111111_1111111111111111_1110110101010101_0001011010100000"; -- -0.07292040437459946
	pesos_i(1236) := b"0000000000000000_0000000000000000_0010100101011110_1111010110000000"; -- 0.16160520911216736
	pesos_i(1237) := b"0000000000000000_0000000000000000_0010101110010000_1100111000000000"; -- 0.17017829418182373
	pesos_i(1238) := b"0000000000000000_0000000000000000_0000100011000110_1110110011110000"; -- 0.03428536280989647
	pesos_i(1239) := b"0000000000000000_0000000000000000_0010011101101101_1101110100000000"; -- 0.15402013063430786
	pesos_i(1240) := b"0000000000000000_0000000000000000_0010111110000010_1101011111000000"; -- 0.1855902522802353
	pesos_i(1241) := b"1111111111111111_1111111111111111_1110010001111111_0000011101100000"; -- -0.10743669420480728
	pesos_i(1242) := b"1111111111111111_1111111111111111_1010000011111011_1011110110000000"; -- -0.37115874886512756
	pesos_i(1243) := b"0000000000000000_0000000000000000_0010000010100100_1010001111000000"; -- 0.12751220166683197
	pesos_i(1244) := b"0000000000000000_0000000000000000_0010111000101110_0011100110000000"; -- 0.18039283156394958
	pesos_i(1245) := b"1111111111111111_1111111111111111_1101101100010010_0010111001000000"; -- -0.14425383508205414
	pesos_i(1246) := b"0000000000000000_0000000000000000_0010111001001101_0011111110000000"; -- 0.18086621165275574
	pesos_i(1247) := b"1111111111111111_1111111111111111_1111001010011111_0101111000010000"; -- -0.052255745977163315
	pesos_i(1248) := b"1111111111111111_1111111111111111_1110100110011101_1101011000000000"; -- -0.08743536472320557
	pesos_i(1249) := b"1111111111111111_1111111111111111_1111010110001100_1000011000000000"; -- -0.0408245325088501
	pesos_i(1250) := b"1111111111111111_1111111111111111_1110010000001100_1111010100100000"; -- -0.10917728394269943
	pesos_i(1251) := b"0000000000000000_0000000000000000_0010001001110101_1000110101000000"; -- 0.13460619747638702
	pesos_i(1252) := b"1111111111111111_1111111111111111_1110001001110000_1000011010000000"; -- -0.11547049880027771
	pesos_i(1253) := b"1111111111111111_1111111111111111_1111001010010001_1101100000110000"; -- -0.05246208980679512
	pesos_i(1254) := b"1111111111111111_1111111111111111_1111001000010001_1011001101100000"; -- -0.054417409002780914
	pesos_i(1255) := b"1111111111111111_1111111111111111_1100011011100001_0010101010000000"; -- -0.22312673926353455
	pesos_i(1256) := b"1111111111111111_1111111111111111_1110111010110100_1011110011100000"; -- -0.06755466014146805
	pesos_i(1257) := b"1111111111111111_1111111111111111_1111111010111100_1000110011000010"; -- -0.0049354578368365765
	pesos_i(1258) := b"1111111111111111_1111111111111111_1111111101111101_1010101010011100"; -- -0.0019887322559952736
	pesos_i(1259) := b"0000000000000000_0000000000000000_0000110100010101_0111111110000000"; -- 0.05110928416252136
	pesos_i(1260) := b"0000000000000000_0000000000000000_0010101110100001_1101010110000000"; -- 0.17043814063072205
	pesos_i(1261) := b"1111111111111111_1111111111111111_1110110100101011_1101100011100000"; -- -0.07354969531297684
	pesos_i(1262) := b"1111111111111111_1111111111111111_1111010101011011_1101011100000000"; -- -0.04156738519668579
	pesos_i(1263) := b"0000000000000000_0000000000000000_0000011000110010_1100000101001000"; -- 0.024211959913372993
	pesos_i(1264) := b"1111111111111111_1111111111111111_1011111001100110_1111001000000000"; -- -0.25624167919158936
	pesos_i(1265) := b"1111111111111111_1111111111111111_1100100101000101_1110100101000000"; -- -0.21377699077129364
	pesos_i(1266) := b"0000000000000000_0000000000000000_0010001010101110_0010011111000000"; -- 0.13546989858150482
	pesos_i(1267) := b"0000000000000000_0000000000000000_0001101001100011_0011101111100000"; -- 0.10307668894529343
	pesos_i(1268) := b"1111111111111111_1111111111111111_1111011101110100_1100100011100000"; -- -0.03337425738573074
	pesos_i(1269) := b"1111111111111111_1111111111111111_1101111001111111_0000101001000000"; -- -0.13087402284145355
	pesos_i(1270) := b"0000000000000000_0000000000000000_0000010001000111_0101010001110000"; -- 0.016713406890630722
	pesos_i(1271) := b"0000000000000000_0000000000000000_0011011101100101_1011010111000000"; -- 0.21639572083950043
	pesos_i(1272) := b"0000000000000000_0000000000000000_0010101111110000_1111110100000000"; -- 0.17164593935012817
	pesos_i(1273) := b"1111111111111111_1111111111111111_1111011101101011_1001111011100000"; -- -0.03351408988237381
	pesos_i(1274) := b"1111111111111111_1111111111111111_1101001110001011_1110000011000000"; -- -0.17364688217639923
	pesos_i(1275) := b"0000000000000000_0000000000000000_0001110100100101_0100010110100000"; -- 0.11384997516870499
	pesos_i(1276) := b"1111111111111111_1111111111111111_1011110101001001_0000101100000000"; -- -0.26060420274734497
	pesos_i(1277) := b"1111111111111111_1111111111111111_1110111101100111_0011101110100000"; -- -0.06483104079961777
	pesos_i(1278) := b"0000000000000000_0000000000000000_0000000101111110_0010101010100010"; -- 0.005831398535519838
	pesos_i(1279) := b"0000000000000000_0000000000000000_0001101010111011_0111111001100000"; -- 0.10442342609167099
	pesos_i(1280) := b"0000000000000000_0000000000000000_0010111100100101_0110101100000000"; -- 0.18416470289230347
	pesos_i(1281) := b"1111111111111111_1111111111111111_1101111100000001_1101100111000000"; -- -0.12887801229953766
	pesos_i(1282) := b"0000000000000000_0000000000000000_0100011100110000_0010011110000000"; -- 0.27807852625846863
	pesos_i(1283) := b"1111111111111111_1111111111111111_1100100111000001_1011000111000000"; -- -0.21188820898532867
	pesos_i(1284) := b"1111111111111111_1111111111111111_0111100111100111_0111000000000000"; -- -0.5238122940063477
	pesos_i(1285) := b"1111111111111111_1111111111111111_0101100111010110_1011000100000000"; -- -0.6490678191184998
	pesos_i(1286) := b"0000000000000000_0000000000000000_0011011010011111_1111011111000000"; -- 0.2133784145116806
	pesos_i(1287) := b"1111111111111111_1111111111111111_1110101111011010_0110011101000000"; -- -0.07869867980480194
	pesos_i(1288) := b"1111111111111111_1111111111111111_1110011101010110_0111010001100000"; -- -0.09633705765008926
	pesos_i(1289) := b"1111111111111111_1111111111111111_1110010100111000_0101011011000000"; -- -0.10460908710956573
	pesos_i(1290) := b"0000000000000000_0000000000000000_0100010110101001_0111001100000000"; -- 0.27211683988571167
	pesos_i(1291) := b"0000000000000000_0000000000000000_0100001001001000_1101100100000000"; -- 0.25892406702041626
	pesos_i(1292) := b"1111111111111111_1111111111111111_1110001000001011_1011010111000000"; -- -0.11700882017612457
	pesos_i(1293) := b"1111111111111111_1111111111111111_1101010001110101_1001001010000000"; -- -0.1700809895992279
	pesos_i(1294) := b"0000000000000000_0000000000000000_0100000111111000_1111110100000000"; -- 0.2577055096626282
	pesos_i(1295) := b"0000000000000000_0000000000000000_0001100110101100_0100010111100000"; -- 0.10028492659330368
	pesos_i(1296) := b"1111111111111111_1111111111111111_1110111011101101_0001101111100000"; -- -0.06669450551271439
	pesos_i(1297) := b"0000000000000000_0000000000000000_0000001000110000_0111111001111000"; -- 0.008552459999918938
	pesos_i(1298) := b"1111111111111111_1111111111111111_0100000100100111_0110101100000000"; -- -0.7454922795295715
	pesos_i(1299) := b"1111111111111111_1111111111111111_1011010100011100_1110011110000000"; -- -0.2925277054309845
	pesos_i(1300) := b"0000000000000000_0000000000000000_0101011011011110_1110110110000000"; -- 0.33933910727500916
	pesos_i(1301) := b"0000000000000000_0000000000000000_0100001000011011_0010101110000000"; -- 0.25822708010673523
	pesos_i(1302) := b"0000000000000000_0000000000000000_0011101110101000_1100101110000000"; -- 0.2330443561077118
	pesos_i(1303) := b"1111111111111111_1111111111111111_1101001111000001_1110001010000000"; -- -0.17282280325889587
	pesos_i(1304) := b"1111111111111111_1111111111111111_1001111111001111_0111001000000000"; -- -0.3757408857345581
	pesos_i(1305) := b"1111111111111111_1111111111111111_1110010111100000_1001001010100000"; -- -0.10204204171895981
	pesos_i(1306) := b"0000000000000000_0000000000000000_0001010100101000_1100001111000000"; -- 0.08265326917171478
	pesos_i(1307) := b"1111111111111111_1111111111111111_1110010101110101_1100001011100000"; -- -0.1036718562245369
	pesos_i(1308) := b"1111111111111111_1111111111111111_1010010111111110_1101101010000000"; -- -0.3515799939632416
	pesos_i(1309) := b"1111111111111111_1111111111111111_1111011111001111_0010111100100000"; -- -0.03199487179517746
	pesos_i(1310) := b"0000000000000000_0000000000000000_0000110000010011_0111111100000000"; -- 0.047172486782073975
	pesos_i(1311) := b"1111111111111111_1111111111111111_1111110101000010_1110111100010000"; -- -0.010697420686483383
	pesos_i(1312) := b"0000000000000000_0000000000000000_0100011101001010_1001001000000000"; -- 0.2784816026687622
	pesos_i(1313) := b"0000000000000000_0000000000000000_0000011100010111_0111111111000000"; -- 0.027702316641807556
	pesos_i(1314) := b"0000000000000000_0000000000000000_0001100111011010_0110100110000000"; -- 0.1009889543056488
	pesos_i(1315) := b"1111111111111111_1111111111111111_1100110100101101_1011100100000000"; -- -0.19852107763290405
	pesos_i(1316) := b"1111111111111111_1111111111111111_0111100111010100_1011010000000000"; -- -0.5240981578826904
	pesos_i(1317) := b"0000000000000000_0000000000000000_0100110111100011_0110011010000000"; -- 0.304251104593277
	pesos_i(1318) := b"0000000000000000_0000000000000000_0000101100100100_1110110000100000"; -- 0.04353214055299759
	pesos_i(1319) := b"0000000000000000_0000000000000000_0010011111100101_1000001011000000"; -- 0.15584580600261688
	pesos_i(1320) := b"1111111111111111_1111111111111111_1011011110000111_0001000010000000"; -- -0.2830953299999237
	pesos_i(1321) := b"1111111111111111_1111111111111111_1010110111001100_1011110100000000"; -- -0.32109469175338745
	pesos_i(1322) := b"1111111111111111_1111111111111111_1111011111001011_1011101000000000"; -- -0.03204762935638428
	pesos_i(1323) := b"1111111111111111_1111111111111111_1011010011011011_0100011010000000"; -- -0.29352912306785583
	pesos_i(1324) := b"0000000000000000_0000000000000000_0000000101111101_1101100111100110"; -- 0.0058265863917768
	pesos_i(1325) := b"0000000000000000_0000000000000000_0100110010010111_0110111110000000"; -- 0.29918572306632996
	pesos_i(1326) := b"1111111111111111_1111111111111111_1000010110100100_1100111010000000"; -- -0.4779540002346039
	pesos_i(1327) := b"1111111111111111_1111111111111111_1111100100011111_0101111010010000"; -- -0.026865091174840927
	pesos_i(1328) := b"1111111111111111_1111111111111111_1100010001101101_0010000101000000"; -- -0.23270981013774872
	pesos_i(1329) := b"0000000000000000_0000000000000000_0011100100101011_1110100100000000"; -- 0.22332626581192017
	pesos_i(1330) := b"0000000000000000_0000000000000000_0000011000111011_0100110001101000"; -- 0.02434232272207737
	pesos_i(1331) := b"0000000000000000_0000000000000000_0001100011111010_0110101000100000"; -- 0.09757102280855179
	pesos_i(1332) := b"1111111111111111_1111111111111111_1111110000011110_0110111100001100"; -- -0.015160617418587208
	pesos_i(1333) := b"1111111111111111_1111111111111111_1111001100101110_1100111001110000"; -- -0.05006704106926918
	pesos_i(1334) := b"0000000000000000_0000000000000000_0010000111011001_0001001001000000"; -- 0.13221849501132965
	pesos_i(1335) := b"0000000000000000_0000000000000000_0001011001111010_0111001101000000"; -- 0.08780594170093536
	pesos_i(1336) := b"1111111111111111_1111111111111111_1011111011110010_0101001010000000"; -- -0.25411495566368103
	pesos_i(1337) := b"0000000000000000_0000000000000000_0101001111101110_0111111110000000"; -- 0.32785794138908386
	pesos_i(1338) := b"1111111111111111_1111111111111111_1110000011001011_0011101111100000"; -- -0.12189889699220657
	pesos_i(1339) := b"0000000000000000_0000000000000000_0100100101100100_0101000010000000"; -- 0.2866869270801544
	pesos_i(1340) := b"0000000000000000_0000000000000000_0010101000100111_0111111100000000"; -- 0.16466516256332397
	pesos_i(1341) := b"1111111111111111_1111111111111111_1001100110000100_1001100000000000"; -- -0.40032052993774414
	pesos_i(1342) := b"0000000000000000_0000000000000000_0101110000011110_0010001000000000"; -- 0.35983479022979736
	pesos_i(1343) := b"0000000000000000_0000000000000000_0010011110101101_1001001011000000"; -- 0.1549922674894333
	pesos_i(1344) := b"1111111111111111_1111111111111111_1011101110010000_1111111110000000"; -- -0.2673187553882599
	pesos_i(1345) := b"1111111111111111_1111111111111111_1110010100101101_0001111010100000"; -- -0.10478027909994125
	pesos_i(1346) := b"1111111111111111_1111111111111111_1111100110001100_1100001111111000"; -- -0.025195838883519173
	pesos_i(1347) := b"0000000000000000_0000000000000000_0001101100000111_1111101111000000"; -- 0.1055905669927597
	pesos_i(1348) := b"0000000000000000_0000000000000000_0010001011010100_1011011000000000"; -- 0.13605821132659912
	pesos_i(1349) := b"0000000000000000_0000000000000000_0011000111000111_1110110100000000"; -- 0.19445687532424927
	pesos_i(1350) := b"1111111111111111_1111111111111111_1100101001001100_0110000101000000"; -- -0.2097720354795456
	pesos_i(1351) := b"1111111111111111_1111111111111111_1101001010110101_1100100010000000"; -- -0.17691370844841003
	pesos_i(1352) := b"0000000000000000_0000000000000000_0101000100011100_1111101010000000"; -- 0.31684842705726624
	pesos_i(1353) := b"0000000000000000_0000000000000000_0000011010100011_0101010101101000"; -- 0.025929773226380348
	pesos_i(1354) := b"1111111111111111_1111111111111111_1111111101011000_0101101110101111"; -- -0.0025580117944628
	pesos_i(1355) := b"0000000000000000_0000000000000000_0001110010101110_1100111000000000"; -- 0.11204230785369873
	pesos_i(1356) := b"1111111111111111_1111111111111111_1011110011011001_1111111110000000"; -- -0.2622986137866974
	pesos_i(1357) := b"0000000000000000_0000000000000000_0001111110010111_0100100011100000"; -- 0.1234021708369255
	pesos_i(1358) := b"1111111111111111_1111111111111111_1100110011100101_1010011100000000"; -- -0.19962078332901
	pesos_i(1359) := b"1111111111111111_1111111111111111_1010111001101000_1110101000000000"; -- -0.31871163845062256
	pesos_i(1360) := b"0000000000000000_0000000000000000_0001011010010000_1011001011100000"; -- 0.0881454274058342
	pesos_i(1361) := b"0000000000000000_0000000000000000_0000011111000010_0010001000101000"; -- 0.03030599094927311
	pesos_i(1362) := b"1111111111111111_1111111111111111_1111101101000101_1101011001111000"; -- -0.018465610221028328
	pesos_i(1363) := b"1111111111111111_1111111111111111_1101011010001111_1101111101000000"; -- -0.1618671864271164
	pesos_i(1364) := b"0000000000000000_0000000000000000_0011101100000010_1000000100000000"; -- 0.23050695657730103
	pesos_i(1365) := b"0000000000000000_0000000000000000_0010010100111110_0000010010000000"; -- 0.1454775631427765
	pesos_i(1366) := b"0000000000000000_0000000000000000_0000011111011001_1101110111011000"; -- 0.03066813014447689
	pesos_i(1367) := b"0000000000000000_0000000000000000_0101010100010110_0101011100000000"; -- 0.33237212896347046
	pesos_i(1368) := b"0000000000000000_0000000000000000_0010000110111000_0010000111000000"; -- 0.13171587884426117
	pesos_i(1369) := b"0000000000000000_0000000000000000_0000111100101110_1011000101010000"; -- 0.059306222945451736
	pesos_i(1370) := b"1111111111111111_1111111111111111_1101011000111110_0110000110000000"; -- -0.1631106436252594
	pesos_i(1371) := b"0000000000000000_0000000000000000_0011011101101110_1010001111000000"; -- 0.21653197705745697
	pesos_i(1372) := b"0000000000000000_0000000000000000_0110000001001010_0100110110000000"; -- 0.3761337697505951
	pesos_i(1373) := b"1111111111111111_1111111111111111_1111000111100111_1010001100000000"; -- -0.05505925416946411
	pesos_i(1374) := b"0000000000000000_0000000000000000_0010101011111011_0001110000000000"; -- 0.1678941249847412
	pesos_i(1375) := b"0000000000000000_0000000000000000_0000001011110011_1001001111110100"; -- 0.011529204435646534
	pesos_i(1376) := b"0000000000000000_0000000000000000_0000101101111000_0001000111010000"; -- 0.04480086639523506
	pesos_i(1377) := b"1111111111111111_1111111111111111_1110110001101010_1101011000000000"; -- -0.07649481296539307
	pesos_i(1378) := b"1111111111111111_1111111111111111_1111000000100111_1010110110010000"; -- -0.06189456209540367
	pesos_i(1379) := b"0000000000000000_0000000000000000_0001000100011001_1010110100100000"; -- 0.06679803878068924
	pesos_i(1380) := b"1111111111111111_1111111111111111_1110110101001110_1011011010100000"; -- -0.0730176791548729
	pesos_i(1381) := b"0000000000000000_0000000000000000_0001011100000110_1010101110100000"; -- 0.08994553238153458
	pesos_i(1382) := b"1111111111111111_1111111111111111_1110000011010011_0011100100100000"; -- -0.1217769905924797
	pesos_i(1383) := b"0000000000000000_0000000000000000_0001110101000010_0110100110100000"; -- 0.1142946258187294
	pesos_i(1384) := b"0000000000000000_0000000000000000_0000010110111010_1110010000110000"; -- 0.022382985800504684
	pesos_i(1385) := b"1111111111111111_1111111111111111_1100100111000000_0110110010000000"; -- -0.21190759539604187
	pesos_i(1386) := b"1111111111111111_1111111111111111_1111101001011000_1111001011101000"; -- -0.022080248221755028
	pesos_i(1387) := b"0000000000000000_0000000000000000_0000100010011110_0100111001100000"; -- 0.03366556018590927
	pesos_i(1388) := b"0000000000000000_0000000000000000_0001111001001111_1001011111100000"; -- 0.11840199679136276
	pesos_i(1389) := b"1111111111111111_1111111111111111_1010111001101110_0110101110000000"; -- -0.31862762570381165
	pesos_i(1390) := b"0000000000000000_0000000000000000_0000111101011001_1111101101100000"; -- 0.059966765344142914
	pesos_i(1391) := b"0000000000000000_0000000000000000_0001011100111001_1101000101000000"; -- 0.09072597324848175
	pesos_i(1392) := b"1111111111111111_1111111111111111_1111111101011000_1111000101100110"; -- -0.002549088094383478
	pesos_i(1393) := b"1111111111111111_1111111111111111_1101000001100010_0000101100000000"; -- -0.18600398302078247
	pesos_i(1394) := b"0000000000000000_0000000000000000_0100010110010010_1101100110000000"; -- 0.27177199721336365
	pesos_i(1395) := b"1111111111111111_1111111111111111_1110001000111011_1100010100000000"; -- -0.11627548933029175
	pesos_i(1396) := b"1111111111111111_1111111111111111_1111111110101010_0101100100100010"; -- -0.001306943129748106
	pesos_i(1397) := b"1111111111111111_1111111111111111_1011000110100101_0001110000000000"; -- -0.3060743808746338
	pesos_i(1398) := b"0000000000000000_0000000000000000_0010001111110011_0100011011000000"; -- 0.14043085277080536
	pesos_i(1399) := b"0000000000000000_0000000000000000_0010111010010011_1111100111000000"; -- 0.18194542825222015
	pesos_i(1400) := b"0000000000000000_0000000000000000_0001001110111110_1010100011000000"; -- 0.07712797820568085
	pesos_i(1401) := b"0000000000000000_0000000000000000_0000111101111001_1010110010110000"; -- 0.06045035645365715
	pesos_i(1402) := b"1111111111111111_1111111111111111_1011101001000111_1110001110000000"; -- -0.2723405659198761
	pesos_i(1403) := b"1111111111111111_1111111111111111_1110001000100100_0010000010000000"; -- -0.1166362464427948
	pesos_i(1404) := b"1111111111111111_1111111111111111_1111101100101011_1010111010101000"; -- -0.018864711746573448
	pesos_i(1405) := b"1111111111111111_1111111111111111_1011111110001110_0111110000000000"; -- -0.25173211097717285
	pesos_i(1406) := b"1111111111111111_1111111111111111_1100010001110000_1101110011000000"; -- -0.23265285789966583
	pesos_i(1407) := b"0000000000000000_0000000000000000_0100110101011010_1001010100000000"; -- 0.30216342210769653
	pesos_i(1408) := b"1111111111111111_1111111111111111_1111101000100001_1000110110010000"; -- -0.022925522178411484
	pesos_i(1409) := b"0000000000000000_0000000000000000_0001100100000011_0010111010100000"; -- 0.09770480543375015
	pesos_i(1410) := b"0000000000000000_0000000000000000_0011100011000000_0110110011000000"; -- 0.22168616950511932
	pesos_i(1411) := b"1111111111111111_1111111111111111_1110100010110111_1000000110100000"; -- -0.09094991534948349
	pesos_i(1412) := b"0000000000000000_0000000000000000_0001100000000001_1011100100000000"; -- 0.09377628564834595
	pesos_i(1413) := b"1111111111111111_1111111111111111_0011111111011000_1101010100000000"; -- -0.7505976557731628
	pesos_i(1414) := b"1111111111111111_1111111111111111_1111100010100010_0011101011111000"; -- -0.0287745613604784
	pesos_i(1415) := b"1111111111111111_1111111111111111_1010010110000011_0101001100000000"; -- -0.35346490144729614
	pesos_i(1416) := b"1111111111111111_1111111111111111_1100101111011001_1010001111000000"; -- -0.20371033251285553
	pesos_i(1417) := b"0000000000000000_0000000000000000_0010100101110101_1011000101000000"; -- 0.16195209324359894
	pesos_i(1418) := b"0000000000000000_0000000000000000_0000011110100010_1010100011001000"; -- 0.029825733974575996
	pesos_i(1419) := b"0000000000000000_0000000000000000_0100001001111110_1011110010000000"; -- 0.25974634289741516
	pesos_i(1420) := b"0000000000000000_0000000000000000_0001111000011010_1001001000100000"; -- 0.1175929382443428
	pesos_i(1421) := b"1111111111111111_1111111111111111_1011111111011101_0011101000000000"; -- -0.2505306005477905
	pesos_i(1422) := b"0000000000000000_0000000000000000_0010000001001011_1001111100000000"; -- 0.1261538863182068
	pesos_i(1423) := b"0000000000000000_0000000000000000_0010011000101011_0001110111000000"; -- 0.14909540116786957
	pesos_i(1424) := b"0000000000000000_0000000000000000_0000010011000111_1001000100100000"; -- 0.01867014914751053
	pesos_i(1425) := b"0000000000000000_0000000000000000_0010011101110011_1110101100000000"; -- 0.15411251783370972
	pesos_i(1426) := b"0000000000000000_0000000000000000_0000010111000000_1010110110111000"; -- 0.022471291944384575
	pesos_i(1427) := b"1111111111111111_1111111111111111_1100100100110011_0100001000000000"; -- -0.21406161785125732
	pesos_i(1428) := b"0000000000000000_0000000000000000_0001010100001001_1101111000100000"; -- 0.08218181878328323
	pesos_i(1429) := b"0000000000000000_0000000000000000_0010000011001001_0001001011000000"; -- 0.12806813418865204
	pesos_i(1430) := b"0000000000000000_0000000000000000_0000001000011110_0100011010010100"; -- 0.008274470455944538
	pesos_i(1431) := b"0000000000000000_0000000000000000_0100101011111000_1110111010000000"; -- 0.29286089539527893
	pesos_i(1432) := b"1111111111111111_1111111111111111_0110001000001010_0011110000000000"; -- -0.6170313358306885
	pesos_i(1433) := b"0000000000000000_0000000000000000_0000110010110010_1001000001000000"; -- 0.04959966242313385
	pesos_i(1434) := b"0000000000000000_0000000000000000_0110100010000000_0011101010000000"; -- 0.40820661187171936
	pesos_i(1435) := b"0000000000000000_0000000000000000_0000100111011111_0000010011110000"; -- 0.03855925425887108
	pesos_i(1436) := b"1111111111111111_1111111111111111_1100111000101000_1100101111000000"; -- -0.19469000399112701
	pesos_i(1437) := b"0000000000000000_0000000000000000_0001101010110010_0010000011100000"; -- 0.10428052395582199
	pesos_i(1438) := b"0000000000000000_0000000000000000_0010010110001000_1010101001000000"; -- 0.146616593003273
	pesos_i(1439) := b"1111111111111111_1111111111111111_1111011000010101_0011011110100000"; -- -0.03873874992132187
	pesos_i(1440) := b"0000000000000000_0000000000000000_0010101000100010_0000111101000000"; -- 0.16458220779895782
	pesos_i(1441) := b"0000000000000000_0000000000000000_0010010100001011_0001001010000000"; -- 0.14470019936561584
	pesos_i(1442) := b"0000000000000000_0000000000000000_0001001010100101_0000101001100000"; -- 0.07283081859350204
	pesos_i(1443) := b"1111111111111111_1111111111111111_1010100100011110_1010101100000000"; -- -0.3393757939338684
	pesos_i(1444) := b"1111111111111111_1111111111111111_1110010000011010_1011011000100000"; -- -0.10896741598844528
	pesos_i(1445) := b"0000000000000000_0000000000000000_0000110010011000_0011101100000000"; -- 0.04919785261154175
	pesos_i(1446) := b"0000000000000000_0000000000000000_0000100110101011_1111100010100000"; -- 0.03778032213449478
	pesos_i(1447) := b"0000000000000000_0000000000000000_0010001000011110_0001010001000000"; -- 0.1332714706659317
	pesos_i(1448) := b"0000000000000000_0000000000000000_0001001100110010_0011101100100000"; -- 0.07498521357774734
	pesos_i(1449) := b"0000000000000000_0000000000000000_0010110100100000_0111010011000000"; -- 0.17627649009227753
	pesos_i(1450) := b"0000000000000000_0000000000000000_0000011101110000_1011001010011000"; -- 0.029063379392027855
	pesos_i(1451) := b"0000000000000000_0000000000000000_0011011101101100_1111101100000000"; -- 0.21650665998458862
	pesos_i(1452) := b"0000000000000000_0000000000000000_0010111001101001_1101111001000000"; -- 0.18130291998386383
	pesos_i(1453) := b"0000000000000000_0000000000000000_0001001101001010_0110111001100000"; -- 0.07535447925329208
	pesos_i(1454) := b"1111111111111111_1111111111111111_1011111110101011_1101010010000000"; -- -0.25128433108329773
	pesos_i(1455) := b"1111111111111111_1111111111111111_1100100011100101_1001011001000000"; -- -0.21524678170681
	pesos_i(1456) := b"0000000000000000_0000000000000000_0011110100100100_0101101011000000"; -- 0.23883597552776337
	pesos_i(1457) := b"1111111111111111_1111111111111111_1110100110100000_1111100000100000"; -- -0.0873875543475151
	pesos_i(1458) := b"1111111111111111_1111111111111111_1101111001001101_1100001011000000"; -- -0.1316259652376175
	pesos_i(1459) := b"0000000000000000_0000000000000000_0101110001110011_0101110010000000"; -- 0.3611352741718292
	pesos_i(1460) := b"0000000000000000_0000000000000000_0010001001101001_1111001000000000"; -- 0.13442909717559814
	pesos_i(1461) := b"1111111111111111_1111111111111111_1101001111000101_0001010001000000"; -- -0.1727740615606308
	pesos_i(1462) := b"1111111111111111_1111111111111111_1111100001111101_1110101000001000"; -- -0.02932870201766491
	pesos_i(1463) := b"0000000000000000_0000000000000000_0010011100001010_1100001111000000"; -- 0.15250800549983978
	pesos_i(1464) := b"1111111111111111_1111111111111111_1111001001101010_1010001110000000"; -- -0.053060322999954224
	pesos_i(1465) := b"0000000000000000_0000000000000000_0111111000111010_0010101110000000"; -- 0.49307510256767273
	pesos_i(1466) := b"0000000000000000_0000000000000000_0000010010010111_0100011100101000"; -- 0.0179333183914423
	pesos_i(1467) := b"0000000000000000_0000000000000000_0010001010111001_0101001010000000"; -- 0.13564029335975647
	pesos_i(1468) := b"0000000000000000_0000000000000000_0010010011011101_0101000100000000"; -- 0.1440020203590393
	pesos_i(1469) := b"0000000000000000_0000000000000000_0001101000010100_1100001110100000"; -- 0.10187933593988419
	pesos_i(1470) := b"1111111111111111_1111111111111111_1101111101001001_0101001111000000"; -- -0.12778736650943756
	pesos_i(1471) := b"0000000000000000_0000000000000000_0010111011100110_1101000000000000"; -- 0.18320941925048828
	pesos_i(1472) := b"1111111111111111_1111111111111111_1111010111010110_0000100000100000"; -- -0.0397028848528862
	pesos_i(1473) := b"0000000000000000_0000000000000000_0010110010110111_1001001000000000"; -- 0.1746760606765747
	pesos_i(1474) := b"0000000000000000_0000000000000000_0001110110111110_1111010110100000"; -- 0.11619506031274796
	pesos_i(1475) := b"0000000000000000_0000000000000000_0010011111101110_0100001111000000"; -- 0.15597938001155853
	pesos_i(1476) := b"1111111111111111_1111111111111111_1111111111111010_1110000111110111"; -- -7.808421651134267e-05
	pesos_i(1477) := b"1111111111111111_1111111111111111_1110101000011110_0111101110100000"; -- -0.08547236770391464
	pesos_i(1478) := b"1111111111111111_1111111111111111_0010110000100011_0101101000000000"; -- -0.8275855779647827
	pesos_i(1479) := b"1111111111111111_1111111111111111_1110000010100011_1000011011000000"; -- -0.12250478565692902
	pesos_i(1480) := b"0000000000000000_0000000000000000_0111001010100110_1110011000000000"; -- 0.44785916805267334
	pesos_i(1481) := b"1111111111111111_1111111111111111_1100100010000100_1111101111000000"; -- -0.2167208343744278
	pesos_i(1482) := b"1111111111111111_1111111111111111_1010101001001000_1110100000000000"; -- -0.3348250389099121
	pesos_i(1483) := b"1111111111111111_1111111111111111_1100110100101111_0111110010000000"; -- -0.19849416613578796
	pesos_i(1484) := b"0000000000000000_0000000000000000_0011111111000000_0010011111000000"; -- 0.24902580678462982
	pesos_i(1485) := b"0000000000000000_0000000000000000_0101101000100110_0111110010000000"; -- 0.35214975476264954
	pesos_i(1486) := b"0000000000000000_0000000000000000_1000100110111000_0000100000000000"; -- 0.5379643440246582
	pesos_i(1487) := b"1111111111111111_1111111111111111_1010111011001100_1101011000000000"; -- -0.31718695163726807
	pesos_i(1488) := b"1111111111111111_1111111111111111_1110011110000010_1000100010100000"; -- -0.09566446393728256
	pesos_i(1489) := b"0000000000000000_0000000000000000_0110011010010001_0001010100000000"; -- 0.4006512761116028
	pesos_i(1490) := b"1111111111111111_1111111111111111_1100111000001101_0011100011000000"; -- -0.1951107531785965
	pesos_i(1491) := b"1111111111111111_1111111111111111_1110100111110101_0011110111000000"; -- -0.08610166609287262
	pesos_i(1492) := b"1111111111111111_1111111111111111_1101001100011000_0000101111000000"; -- -0.1754143387079239
	pesos_i(1493) := b"0000000000000000_0000000000000000_0000100110100000_1110110011100000"; -- 0.03761177510023117
	pesos_i(1494) := b"1111111111111111_1111111111111111_1111110100000010_1011001100010100"; -- -0.011677558533847332
	pesos_i(1495) := b"1111111111111111_1111111111111111_1100100100010011_1000000010000000"; -- -0.21454617381095886
	pesos_i(1496) := b"0000000000000000_0000000000000000_0010011110010110_0010000011000000"; -- 0.1546345204114914
	pesos_i(1497) := b"1111111111111111_1111111111111111_1111100110100111_1110100101100000"; -- -0.024781621992588043
	pesos_i(1498) := b"0000000000000000_0000000000000000_0010011011111010_0100000000000000"; -- 0.15225601196289062
	pesos_i(1499) := b"1111111111111111_1111111111111111_1111110100000100_1010110011010100"; -- -0.011647413484752178
	pesos_i(1500) := b"0000000000000000_0000000000000000_0001011100011001_1000101100000000"; -- 0.09023350477218628
	pesos_i(1501) := b"0000000000000000_0000000000000000_0001101111000110_0011010100100000"; -- 0.10849315673112869
	pesos_i(1502) := b"0000000000000000_0000000000000000_0100110011111100_0001000100000000"; -- 0.3007212281227112
	pesos_i(1503) := b"1111111111111111_1111111111111111_1100111100101011_0011100100000000"; -- -0.1907467246055603
	pesos_i(1504) := b"0000000000000000_0000000000000000_0100101001001010_0110101010000000"; -- 0.2901979982852936
	pesos_i(1505) := b"1111111111111111_1111111111111111_1110101000100100_0110110110000000"; -- -0.0853816568851471
	pesos_i(1506) := b"1111111111111111_1111111111111111_1111010000011110_1001001000100000"; -- -0.046408526599407196
	pesos_i(1507) := b"0000000000000000_0000000000000000_0010011010110111_1100101100000000"; -- 0.1512419581413269
	pesos_i(1508) := b"0000000000000000_0000000000000000_0001101001100100_1100011100100000"; -- 0.1031002476811409
	pesos_i(1509) := b"0000000000000000_0000000000000000_0011001101010000_0111100110000000"; -- 0.2004466950893402
	pesos_i(1510) := b"1111111111111111_1111111111111111_1111000100100101_1001100101010000"; -- -0.05802003666758537
	pesos_i(1511) := b"0000000000000000_0000000000000000_0100110101001100_0001111100000000"; -- 0.30194276571273804
	pesos_i(1512) := b"1111111111111111_1111111111111111_1110110001111001_0000110000000000"; -- -0.0762779712677002
	pesos_i(1513) := b"1111111111111111_1111111111111111_1001010101111101_0010010000000000"; -- -0.4160592555999756
	pesos_i(1514) := b"0000000000000000_0000000000000000_0100010100010000_0110100010000000"; -- 0.26978161931037903
	pesos_i(1515) := b"0000000000000000_0000000000000000_0010000011111101_1010011110000000"; -- 0.12887045741081238
	pesos_i(1516) := b"1111111111111111_1111111111111111_1011110000111000_1011111000000000"; -- -0.2647591829299927
	pesos_i(1517) := b"1111111111111111_1111111111111111_1111001011000110_1110010010100000"; -- -0.051652632653713226
	pesos_i(1518) := b"0000000000000000_0000000000000000_0000111100001001_1001101111100000"; -- 0.058740369975566864
	pesos_i(1519) := b"0000000000000000_0000000000000000_0001101001000001_0011000110000000"; -- 0.10255727171897888
	pesos_i(1520) := b"0000000000000000_0000000000000000_0000011011110100_0101010110111000"; -- 0.02716575376689434
	pesos_i(1521) := b"1111111111111111_1111111111111111_1101110011011011_0011000111000000"; -- -0.13728035986423492
	pesos_i(1522) := b"1111111111111111_1111111111111111_1100011011010001_1011001001000000"; -- -0.2233627885580063
	pesos_i(1523) := b"1111111111111111_1111111111111111_1000111011000111_0001111000000000"; -- -0.44227421283721924
	pesos_i(1524) := b"1111111111111111_1111111111111111_1100000100000100_1000110010000000"; -- -0.24602434039115906
	pesos_i(1525) := b"1111111111111111_1111111111111111_1111110001101100_1001000110100100"; -- -0.013968369923532009
	pesos_i(1526) := b"1111111111111111_1111111111111111_1101101010110011_1110101100000000"; -- -0.14569216966629028
	pesos_i(1527) := b"0000000000000000_0000000000000000_0100101110111110_1111010110000000"; -- 0.29588255286216736
	pesos_i(1528) := b"1111111111111111_1111111111111111_1100000101111101_1010101000000000"; -- -0.24417626857757568
	pesos_i(1529) := b"1111111111111111_1111111111111111_1111101111100101_1111110000010000"; -- -0.016021963208913803
	pesos_i(1530) := b"1111111111111111_1111111111111111_1110011110111001_0100001110100000"; -- -0.09482934325933456
	pesos_i(1531) := b"1111111111111111_1111111111111111_1111001111010000_0010000101000000"; -- -0.04760544002056122
	pesos_i(1532) := b"1111111111111111_1111111111111111_1101001100101100_1011000100000000"; -- -0.17509931325912476
	pesos_i(1533) := b"0000000000000000_0000000000000000_0010100000010010_0101000111000000"; -- 0.1565295308828354
	pesos_i(1534) := b"0000000000000000_0000000000000000_0000011011000011_0111100101111000"; -- 0.02642020396888256
	pesos_i(1535) := b"0000000000000000_0000000000000000_0110101011010010_1011001110000000"; -- 0.4172775447368622
	pesos_i(1536) := b"1111111111111111_1111111111111111_1111001011000111_0001011111100000"; -- -0.05164957791566849
	pesos_i(1537) := b"1111111111111111_1111111111111111_1101001110000111_1101011001000000"; -- -0.17370854318141937
	pesos_i(1538) := b"0000000000000000_0000000000000000_0001100110000101_0011111100100000"; -- 0.09968943148851395
	pesos_i(1539) := b"1111111111111111_1111111111111111_1101011000111000_0001010010000000"; -- -0.1632067859172821
	pesos_i(1540) := b"0000000000000000_0000000000000000_0010110100110110_1010010110000000"; -- 0.17661508917808533
	pesos_i(1541) := b"1111111111111111_1111111111111111_0101011111000000_0001110100000000"; -- -0.6572248339653015
	pesos_i(1542) := b"0000000000000000_0000000000000000_0100110101011001_1111000110000000"; -- 0.30215367674827576
	pesos_i(1543) := b"1111111111111111_1111111111111111_1110001110110011_1100101001000000"; -- -0.11053787171840668
	pesos_i(1544) := b"1111111111111111_1111111111111111_1011010000000010_0001010010000000"; -- -0.2968432605266571
	pesos_i(1545) := b"0000000000000000_0000000000000000_0100111001000001_1010100010000000"; -- 0.30568936467170715
	pesos_i(1546) := b"1111111111111111_1111111111111111_1100010101001111_0110110111000000"; -- -0.2292567640542984
	pesos_i(1547) := b"1111111111111111_1111111111111111_1101101110000101_0110110011000000"; -- -0.14249534904956818
	pesos_i(1548) := b"0000000000000000_0000000000000000_0011101101000010_0011000011000000"; -- 0.2314787358045578
	pesos_i(1549) := b"1111111111111111_1111111111111111_1001101011011010_1111011100000000"; -- -0.3950963616371155
	pesos_i(1550) := b"1111111111111111_1111111111111111_1111010111111111_0000001101100000"; -- -0.03907755762338638
	pesos_i(1551) := b"1111111111111111_1111111111111111_1110000010001110_0011110011000000"; -- -0.1228296309709549
	pesos_i(1552) := b"0000000000000000_0000000000000000_0010001010110010_0101000011000000"; -- 0.1355333775281906
	pesos_i(1553) := b"0000000000000000_0000000000000000_0101110001111000_1000100100000000"; -- 0.36121422052383423
	pesos_i(1554) := b"0000000000000000_0000000000000000_0110100001001110_1010100010000000"; -- 0.40745022892951965
	pesos_i(1555) := b"0000000000000000_0000000000000000_0100010000000111_0111101010000000"; -- 0.2657391130924225
	pesos_i(1556) := b"0000000000000000_0000000000000000_0100011010111001_1010111100000000"; -- 0.2762708067893982
	pesos_i(1557) := b"0000000000000000_0000000000000000_0011011110011111_1001110111000000"; -- 0.21727930009365082
	pesos_i(1558) := b"0000000000000000_0000000000000000_0010100100101111_0110111011000000"; -- 0.16088001430034637
	pesos_i(1559) := b"0000000000000000_0000000000000000_0001100011100010_0001000101100000"; -- 0.09719952195882797
	pesos_i(1560) := b"1111111111111111_1111111111111111_0110100010100000_0010010000000000"; -- -0.5913064479827881
	pesos_i(1561) := b"1111111111111111_1111111111111111_1011110000000101_1000100110000000"; -- -0.2655405104160309
	pesos_i(1562) := b"0000000000000000_0000000000000000_0010110110010100_0101101011000000"; -- 0.17804495990276337
	pesos_i(1563) := b"0000000000000000_0000000000000000_0101111010011110_1110101100000000"; -- 0.3696123957633972
	pesos_i(1564) := b"1111111111111111_1111111111111111_0110111110101011_1111111100000000"; -- -0.5637817978858948
	pesos_i(1565) := b"0000000000000000_0000000000000000_0011100110000110_0100110000000000"; -- 0.22470545768737793
	pesos_i(1566) := b"0000000000000000_0000000000000000_0011001001100101_0000001101000000"; -- 0.19685383141040802
	pesos_i(1567) := b"0000000000000000_0000000000000000_0001000010000011_0110011110000000"; -- 0.06450507044792175
	pesos_i(1568) := b"1111111111111111_1111111111111111_0100111110011111_0100011100000000"; -- -0.6889758706092834
	pesos_i(1569) := b"0000000000000000_0000000000000000_0011100000111110_1010110001000000"; -- 0.21970631182193756
	pesos_i(1570) := b"0000000000000000_0000000000000000_0011001110100110_0100000101000000"; -- 0.2017555981874466
	pesos_i(1571) := b"1111111111111111_1111111111111111_1011010101001001_1100010100000000"; -- -0.29184311628341675
	pesos_i(1572) := b"0000000000000000_0000000000000000_0000101100001001_0100011100000000"; -- 0.04311031103134155
	pesos_i(1573) := b"0000000000000000_0000000000000000_0000000011110011_1101001100000001"; -- 0.003720462555065751
	pesos_i(1574) := b"1111111111111111_1111111111111111_1111100111100000_0100110010110000"; -- -0.023921210318803787
	pesos_i(1575) := b"0000000000000000_0000000000000000_0011010001100011_0001101110000000"; -- 0.20463725924491882
	pesos_i(1576) := b"0000000000000000_0000000000000000_0111000111001001_0111011100000000"; -- 0.44448035955429077
	pesos_i(1577) := b"0000000000000000_0000000000000000_0100111111011010_1101100010000000"; -- 0.31193307042121887
	pesos_i(1578) := b"0000000000000000_0000000000000000_0001100000100100_1100000110100000"; -- 0.09431085735559464
	pesos_i(1579) := b"0000000000000000_0000000000000000_0010000001101110_0100000011000000"; -- 0.1266823261976242
	pesos_i(1580) := b"1111111111111111_1111111111111111_1101100000001101_1101111001000000"; -- -0.15603838860988617
	pesos_i(1581) := b"0000000000000000_0000000000000000_0011010100011100_1100011010000000"; -- 0.20747032761573792
	pesos_i(1582) := b"1111111111111111_1111111111111111_1110011010101011_1110001010000000"; -- -0.09893974661827087
	pesos_i(1583) := b"1111111111111111_1111111111111111_1110100100100101_1101011001000000"; -- -0.08926640450954437
	pesos_i(1584) := b"0000000000000000_0000000000000000_1000010110110111_0000011000000000"; -- 0.5223239660263062
	pesos_i(1585) := b"1111111111111111_1111111111111111_1101010101101000_0100001011000000"; -- -0.16637785732746124
	pesos_i(1586) := b"1111111111111111_1111111111111111_1011111010111110_0100110000000000"; -- -0.25490880012512207
	pesos_i(1587) := b"0000000000000000_0000000000000000_0110011100000111_1011100100000000"; -- 0.40246158838272095
	pesos_i(1588) := b"0000000000000000_0000000000000000_0011010100000110_1011001101000000"; -- 0.207133486866951
	pesos_i(1589) := b"1111111111111111_1111111111111111_1110000111111110_0011010100100000"; -- -0.11721485108137131
	pesos_i(1590) := b"0000000000000000_0000000000000000_0100100111100000_0101011010000000"; -- 0.28857937455177307
	pesos_i(1591) := b"0000000000000000_0000000000000000_0011001001100010_0010110000000000"; -- 0.19681048393249512
	pesos_i(1592) := b"1111111111111111_1111111111111111_1110110110100001_1010111011100000"; -- -0.0717516615986824
	pesos_i(1593) := b"0000000000000000_0000000000000000_0001000110011100_0001101100000000"; -- 0.06878823041915894
	pesos_i(1594) := b"1111111111111111_1111111111111111_1101111100111001_0111101100000000"; -- -0.12802916765213013
	pesos_i(1595) := b"0000000000000000_0000000000000000_0010110001011111_0100101000000000"; -- 0.17332899570465088
	pesos_i(1596) := b"0000000000000000_0000000000000000_0010011100001010_0010001000000000"; -- 0.15249836444854736
	pesos_i(1597) := b"0000000000000000_0000000000000000_0100100001100000_0001110010000000"; -- 0.2827165424823761
	pesos_i(1598) := b"1111111111111111_1111111111111111_1001000011100011_0010110000000000"; -- -0.4340336322784424
	pesos_i(1599) := b"0000000000000000_0000000000000000_0100110011001001_1011101100000000"; -- 0.2999531626701355
	pesos_i(1600) := b"1111111111111111_1111111111111111_1100111110001100_1101100011000000"; -- -0.18925710022449493
	pesos_i(1601) := b"1111111111111111_1111111111111111_1000101101111100_1111001100000000"; -- -0.4551246762275696
	pesos_i(1602) := b"0000000000000000_0000000000000000_0100101010010001_1001000000000000"; -- 0.29128360748291016
	pesos_i(1603) := b"0000000000000000_0000000000000000_0111011111010011_0111110110000000"; -- 0.4680708348751068
	pesos_i(1604) := b"1111111111111111_1111111111111111_1001011111010101_1100110000000000"; -- -0.4068939685821533
	pesos_i(1605) := b"0000000000000000_0000000000000000_0010000001011100_0101010111000000"; -- 0.1264089196920395
	pesos_i(1606) := b"1111111111111111_1111111111111111_0111111010000011_0100010100000000"; -- -0.505809485912323
	pesos_i(1607) := b"0000000000000000_0000000000000000_0001110001110010_0100100110000000"; -- 0.11111888289451599
	pesos_i(1608) := b"1111111111111111_1111111111111111_1111111010000001_0111100101010100"; -- -0.005836884491145611
	pesos_i(1609) := b"1111111111111111_1111111111111111_1110010100111110_0111010001100000"; -- -0.10451576858758926
	pesos_i(1610) := b"1111111111111111_1111111111111111_1100011000000010_1101110110000000"; -- -0.22651877999305725
	pesos_i(1611) := b"1111111111111111_1111111111111111_1111000010000100_0000100101110000"; -- -0.06048527732491493
	pesos_i(1612) := b"0000000000000000_0000000000000000_0111011100110111_1010111010000000"; -- 0.4656933844089508
	pesos_i(1613) := b"0000000000000000_0000000000000000_0101000000010100_0111000010000000"; -- 0.31281188130378723
	pesos_i(1614) := b"0000000000000000_0000000000000000_0010011001100110_0110000101000000"; -- 0.1499996930360794
	pesos_i(1615) := b"1111111111111111_1111111111111111_1111110101111000_1011100010011100"; -- -0.009876691736280918
	pesos_i(1616) := b"1111111111111111_1111111111111111_1101110111110001_1100101010000000"; -- -0.13302931189537048
	pesos_i(1617) := b"0000000000000000_0000000000000000_0011101010110011_0110011100000000"; -- 0.22929996252059937
	pesos_i(1618) := b"1111111111111111_1111111111111111_1111000100111100_1101100001000000"; -- -0.05766533315181732
	pesos_i(1619) := b"1111111111111111_1111111111111111_1110000011100111_1111011000000000"; -- -0.12146055698394775
	pesos_i(1620) := b"1111111111111111_1111111111111111_1010111001101110_0111010000000000"; -- -0.31862711906433105
	pesos_i(1621) := b"1111111111111111_1111111111111111_1101110010101110_1101110101000000"; -- -0.13795678317546844
	pesos_i(1622) := b"0000000000000000_0000000000000000_0010010000011100_1011010110000000"; -- 0.14106306433677673
	pesos_i(1623) := b"1111111111111111_1111111111111111_0110100000001111_0011101000000000"; -- -0.5935176610946655
	pesos_i(1624) := b"0000000000000000_0000000000000000_0010110100101110_1001111100000000"; -- 0.1764926314353943
	pesos_i(1625) := b"1111111111111111_1111111111111111_1110010100110011_1010101001100000"; -- -0.10468039661645889
	pesos_i(1626) := b"0000000000000000_0000000000000000_0010110011011001_0111011100000000"; -- 0.17519325017929077
	pesos_i(1627) := b"1111111111111111_1111111111111111_1101100000100101_1110000100000000"; -- -0.15567201375961304
	pesos_i(1628) := b"1111111111111111_1111111111111111_1011001110101000_0110101010000000"; -- -0.2982114255428314
	pesos_i(1629) := b"0000000000000000_0000000000000000_0011010000001001_0100110011000000"; -- 0.203266903758049
	pesos_i(1630) := b"0000000000000000_0000000000000000_0000000010010111_1111110000110000"; -- 0.002319108694791794
	pesos_i(1631) := b"0000000000000000_0000000000000000_0011100111001111_1100001110000000"; -- 0.2258264720439911
	pesos_i(1632) := b"0000000000000000_0000000000000000_0011001100000101_0110111000000000"; -- 0.1993016004562378
	pesos_i(1633) := b"1111111111111111_1111111111111111_1111001100001100_0010001100100000"; -- -0.050596050918102264
	pesos_i(1634) := b"0000000000000000_0000000000000000_0110001000001110_0000101100000000"; -- 0.38302677869796753
	pesos_i(1635) := b"0000000000000000_0000000000000000_0011101000101101_1100101011000000"; -- 0.2272612303495407
	pesos_i(1636) := b"0000000000000000_0000000000000000_0001111100010100_0110111100100000"; -- 0.12140554934740067
	pesos_i(1637) := b"0000000000000000_0000000000000000_0011101010001101_1100011100000000"; -- 0.2287258505821228
	pesos_i(1638) := b"1111111111111111_1111111111111111_1010101001100100_1101001110000000"; -- -0.33439901471138
	pesos_i(1639) := b"0000000000000000_0000000000000000_0111010001000110_0001110000000000"; -- 0.4541947841644287
	pesos_i(1640) := b"0000000000000000_0000000000000000_0010001010001100_1111011100000000"; -- 0.13496345281600952
	pesos_i(1641) := b"1111111111111111_1111111111111111_1011011000111111_0001010000000000"; -- -0.288100004196167
	pesos_i(1642) := b"0000000000000000_0000000000000000_0010111110000111_1001100110000000"; -- 0.18566283583641052
	pesos_i(1643) := b"0000000000000000_0000000000000000_0001001100100010_0110110111000000"; -- 0.0747440904378891
	pesos_i(1644) := b"0000000000000000_0000000000000000_0011100111010001_1001100110000000"; -- 0.22585448622703552
	pesos_i(1645) := b"1111111111111111_1111111111111111_1110000011110011_0001101010000000"; -- -0.12129053473472595
	pesos_i(1646) := b"0000000000000000_0000000000000000_0011010000110111_1000100111000000"; -- 0.2039724439382553
	pesos_i(1647) := b"0000000000000000_0000000000000000_0010100101110101_0010100100000000"; -- 0.1619439721107483
	pesos_i(1648) := b"0000000000000000_0000000000000000_0000000100111011_0000101010010100"; -- 0.004807149060070515
	pesos_i(1649) := b"1111111111111111_1111111111111111_1101000110111100_1111110001000000"; -- -0.1807100623846054
	pesos_i(1650) := b"1111111111111111_1111111111111111_1111110101101110_1010010011100000"; -- -0.010030455887317657
	pesos_i(1651) := b"1111111111111111_1111111111111111_1001010011010011_1010010000000000"; -- -0.41864562034606934
	pesos_i(1652) := b"0000000000000000_0000000000000000_0000000110110001_1110101001000110"; -- 0.006621019449084997
	pesos_i(1653) := b"0000000000000000_0000000000000000_0100000100000110_1001000010000000"; -- 0.25400641560554504
	pesos_i(1654) := b"1111111111111111_1111111111111111_1110100101100110_0101110001100000"; -- -0.08828184753656387
	pesos_i(1655) := b"0000000000000000_0000000000000000_0100110010100100_1011000010000000"; -- 0.29938796162605286
	pesos_i(1656) := b"1111111111111111_1111111111111111_1010001011111101_1001001100000000"; -- -0.3633182644844055
	pesos_i(1657) := b"0000000000000000_0000000000000000_0001001110011001_1110010000000000"; -- 0.07656693458557129
	pesos_i(1658) := b"0000000000000000_0000000000000000_0010011111011000_0110000101000000"; -- 0.1556454449892044
	pesos_i(1659) := b"1111111111111111_1111111111111111_1101111010100011_1110011000000000"; -- -0.13031160831451416
	pesos_i(1660) := b"0000000000000000_0000000000000000_0010110101101001_1111101100000000"; -- 0.17739838361740112
	pesos_i(1661) := b"0000000000000000_0000000000000000_0001100101001000_1111001101000000"; -- 0.09876938164234161
	pesos_i(1662) := b"0000000000000000_0000000000000000_0010100000000010_0000001001000000"; -- 0.15628065168857574
	pesos_i(1663) := b"0000000000000000_0000000000000000_1010111101010101_1101110100000000"; -- 0.6849039196968079
	pesos_i(1664) := b"1111111111111111_1111111111111111_1111100101010001_1000001001100000"; -- -0.02610001713037491
	pesos_i(1665) := b"1111111111111111_1111111111111111_1111111001000111_0001110011000000"; -- -0.0067274123430252075
	pesos_i(1666) := b"0000000000000000_0000000000000000_0000100000111001_1011110010100000"; -- 0.03213099390268326
	pesos_i(1667) := b"0000000000000000_0000000000000000_0011011000111111_0111001111000000"; -- 0.21190570294857025
	pesos_i(1668) := b"0000000000000000_0000000000000000_0100101010011110_1100000000000000"; -- 0.2914848327636719
	pesos_i(1669) := b"1111111111111111_1111111111111111_0101001110100101_1101000000000000"; -- -0.6732511520385742
	pesos_i(1670) := b"0000000000000000_0000000000000000_0010010010110111_1000100111000000"; -- 0.1434255689382553
	pesos_i(1671) := b"0000000000000000_0000000000000000_0001100110100010_1011011010100000"; -- 0.1001390591263771
	pesos_i(1672) := b"0000000000000000_0000000000000000_0011100100010000_0100100001000000"; -- 0.22290469706058502
	pesos_i(1673) := b"0000000000000000_0000000000000000_0000100100010010_1011100011000000"; -- 0.03544192016124725
	pesos_i(1674) := b"0000000000000000_0000000000000000_0011010100010011_1101000100000000"; -- 0.20733362436294556
	pesos_i(1675) := b"1111111111111111_1111111111111111_0101011011111101_0111001100000000"; -- -0.6601951718330383
	pesos_i(1676) := b"0000000000000000_0000000000000000_0001000000001001_1111010100000000"; -- 0.06265193223953247
	pesos_i(1677) := b"0000000000000000_0000000000000000_0001011001001111_0010011000100000"; -- 0.08714521676301956
	pesos_i(1678) := b"0000000000000000_0000000000000000_0000110001001110_1000110001010000"; -- 0.04807354882359505
	pesos_i(1679) := b"1111111111111111_1111111111111111_1111100011111011_0001101101101000"; -- -0.027418410405516624
	pesos_i(1680) := b"0000000000000000_0000000000000000_0001101010000100_1110000100000000"; -- 0.10359007120132446
	pesos_i(1681) := b"0000000000000000_0000000000000000_0010010000100111_0110011010000000"; -- 0.14122620224952698
	pesos_i(1682) := b"0000000000000000_0000000000000000_0011000001110110_1011101110000000"; -- 0.18931171298027039
	pesos_i(1683) := b"0000000000000000_0000000000000000_0001111100111111_0010010110000000"; -- 0.12205728888511658
	pesos_i(1684) := b"0000000000000000_0000000000000000_0001001111000110_0101110100100000"; -- 0.07724554091691971
	pesos_i(1685) := b"1111111111111111_1111111111111111_1111000101001110_0011101000000000"; -- -0.05740010738372803
	pesos_i(1686) := b"0000000000000000_0000000000000000_0000010111001101_0101010000100000"; -- 0.02266431599855423
	pesos_i(1687) := b"1111111111111111_1111111111111111_1111011110110000_1111111011010000"; -- -0.03245551511645317
	pesos_i(1688) := b"1111111111111111_1111111111111111_1101001100000111_0010011101000000"; -- -0.17567209899425507
	pesos_i(1689) := b"0000000000000000_0000000000000000_0010100100010101_0111110010000000"; -- 0.16048410534858704
	pesos_i(1690) := b"0000000000000000_0000000000000000_0000100101110111_1001111101110000"; -- 0.036981549113988876
	pesos_i(1691) := b"1111111111111111_1111111111111111_1111011001001000_0111100011010000"; -- -0.03795666620135307
	pesos_i(1692) := b"1111111111111111_1111111111111111_0011011110101100_0111010000000000"; -- -0.782524824142456
	pesos_i(1693) := b"0000000000000000_0000000000000000_0001110010101000_1011110111000000"; -- 0.11194978654384613
	pesos_i(1694) := b"1111111111111111_1111111111111111_1100011010101001_0101001000000000"; -- -0.22397887706756592
	pesos_i(1695) := b"0000000000000000_0000000000000000_0000111110101100_0000100101010000"; -- 0.06121881678700447
	pesos_i(1696) := b"1111111111111111_1111111111111111_0101011101100111_0011000100000000"; -- -0.6585816740989685
	pesos_i(1697) := b"0000000000000000_0000000000000000_0101010111110010_0011001010000000"; -- 0.33572688698768616
	pesos_i(1698) := b"0000000000000000_0000000000000000_0010000011111011_1100001101000000"; -- 0.1288415938615799
	pesos_i(1699) := b"0000000000000000_0000000000000000_0000111010110010_1111100111110000"; -- 0.05741846188902855
	pesos_i(1700) := b"0000000000000000_0000000000000000_0010011100010111_0111001111000000"; -- 0.15270160138607025
	pesos_i(1701) := b"0000000000000000_0000000000000000_0001111011110011_1000100000100000"; -- 0.12090349942445755
	pesos_i(1702) := b"0000000000000000_0000000000000000_0010011011011111_1000000110000000"; -- 0.1518479287624359
	pesos_i(1703) := b"1111111111111111_1111111111111111_1101001011100111_1110101110000000"; -- -0.1761486828327179
	pesos_i(1704) := b"0000000000000000_0000000000000000_0110010100101100_1110100100000000"; -- 0.39521652460098267
	pesos_i(1705) := b"0000000000000000_0000000000000000_0000110011001101_1001010010110000"; -- 0.05001191422343254
	pesos_i(1706) := b"1111111111111111_1111111111111111_1101001010011000_0011000001000000"; -- -0.1773652881383896
	pesos_i(1707) := b"1111111111111111_1111111111111111_1111011000000001_0110010111010000"; -- -0.039041172713041306
	pesos_i(1708) := b"1111111111111111_1111111111111111_1100000011011011_0010110111000000"; -- -0.24665559828281403
	pesos_i(1709) := b"0000000000000000_0000000000000000_0001111000000010_1111111100000000"; -- 0.11723321676254272
	pesos_i(1710) := b"0000000000000000_0000000000000000_0000000110010011_1000101101110110"; -- 0.0061576045118272305
	pesos_i(1711) := b"0000000000000000_0000000000000000_0011000010100100_0001000110000000"; -- 0.19000348448753357
	pesos_i(1712) := b"0000000000000000_0000000000000000_0011100000000011_0101111010000000"; -- 0.21880140900611877
	pesos_i(1713) := b"0000000000000000_0000000000000000_0010011110010001_0100000101000000"; -- 0.1545601636171341
	pesos_i(1714) := b"0000000000000000_0000000000000000_0011000111110111_1011110110000000"; -- 0.19518646597862244
	pesos_i(1715) := b"0000000000000000_0000000000000000_0100101110011011_0100000100000000"; -- 0.2953377366065979
	pesos_i(1716) := b"1111111111111111_1111111111111111_1111110101011110_0001100111000000"; -- -0.010282889008522034
	pesos_i(1717) := b"0000000000000000_0000000000000000_0000111110100101_1001000110110000"; -- 0.061120133846998215
	pesos_i(1718) := b"0000000000000000_0000000000000000_0000110101010111_0100101111100000"; -- 0.05211328715085983
	pesos_i(1719) := b"1111111111111111_1111111111111111_1111110100011011_1110110000010100"; -- -0.011292691342532635
	pesos_i(1720) := b"0000000000000000_0000000000000000_0101010001110111_0011001010000000"; -- 0.32994380593299866
	pesos_i(1721) := b"1111111111111111_1111111111111111_1101000101000010_1010110111000000"; -- -0.18257631361484528
	pesos_i(1722) := b"1111111111111111_1111111111111111_1110100001011101_0100000010000000"; -- -0.09232708811759949
	pesos_i(1723) := b"1111111111111111_1111111111111111_1111001101001100_0000001101100000"; -- -0.04962138086557388
	pesos_i(1724) := b"0000000000000000_0000000000000000_0010010101000001_0110011001000000"; -- 0.14552916586399078
	pesos_i(1725) := b"0000000000000000_0000000000000000_0011000000011101_1001001110000000"; -- 0.18795129656791687
	pesos_i(1726) := b"1111111111111111_1111111111111111_1101111110100001_0110111001000000"; -- -0.126443013548851
	pesos_i(1727) := b"0000000000000000_0000000000000000_0010001110110110_0011100000000000"; -- 0.13949918746948242
	pesos_i(1728) := b"0000000000000000_0000000000000000_0000001111001011_1101101110110000"; -- 0.014829378575086594
	pesos_i(1729) := b"1111111111111111_1111111111111111_1010110101110100_1110111000000000"; -- -0.32243454456329346
	pesos_i(1730) := b"1111111111111111_1111111111111111_1111001110010101_1111101110000000"; -- -0.04849269986152649
	pesos_i(1731) := b"0000000000000000_0000000000000000_0011000000000110_1110001110000000"; -- 0.1876051127910614
	pesos_i(1732) := b"0000000000000000_0000000000000000_0001011100011100_1001000110000000"; -- 0.09027966856956482
	pesos_i(1733) := b"0000000000000000_0000000000000000_0001011010110001_1010000010000000"; -- 0.08864787220954895
	pesos_i(1734) := b"1111111111111111_1111111111111111_1111000111001000_0011101101010000"; -- -0.05553845688700676
	pesos_i(1735) := b"0000000000000000_0000000000000000_0011101011100101_1001010100000000"; -- 0.23006564378738403
	pesos_i(1736) := b"0000000000000000_0000000000000000_0000001111011011_1100110010101000"; -- 0.015072623267769814
	pesos_i(1737) := b"0000000000000000_0000000000000000_0001000001110011_0111111110100000"; -- 0.06426236778497696
	pesos_i(1738) := b"0000000000000000_0000000000000000_0010001111000001_1111010011000000"; -- 0.13967828452587128
	pesos_i(1739) := b"1111111111111111_1111111111111111_1110111011101101_0011000011100000"; -- -0.0666932538151741
	pesos_i(1740) := b"0000000000000000_0000000000000000_0101001110111101_0011001100000000"; -- 0.32710570096969604
	pesos_i(1741) := b"0000000000000000_0000000000000000_0001010100011110_0110111111000000"; -- 0.08249567449092865
	pesos_i(1742) := b"1111111111111111_1111111111111111_1100010111111111_0000111100000000"; -- -0.22657686471939087
	pesos_i(1743) := b"0000000000000000_0000000000000000_0110010000010110_0100000010000000"; -- 0.390964537858963
	pesos_i(1744) := b"1111111111111111_1111111111111111_1110111101111101_0111001101000000"; -- -0.06449203193187714
	pesos_i(1745) := b"0000000000000000_0000000000000000_0101010011111011_0101101100000000"; -- 0.33196038007736206
	pesos_i(1746) := b"0000000000000000_0000000000000000_0000010011101111_1010000000010000"; -- 0.01928139105439186
	pesos_i(1747) := b"0000000000000000_0000000000000000_0100111110011110_0011100110000000"; -- 0.3110080659389496
	pesos_i(1748) := b"0000000000000000_0000000000000000_0010101011100100_1000010101000000"; -- 0.16754944622516632
	pesos_i(1749) := b"0000000000000000_0000000000000000_0010100011011010_1001101110000000"; -- 0.15958568453788757
	pesos_i(1750) := b"0000000000000000_0000000000000000_0000110011101111_1000000000010000"; -- 0.05052948370575905
	pesos_i(1751) := b"1111111111111111_1111111111111111_1011010101010000_1011011000000000"; -- -0.2917371988296509
	pesos_i(1752) := b"0000000000000000_0000000000000000_0000101001001111_1011010010010000"; -- 0.040278706699609756
	pesos_i(1753) := b"0000000000000000_0000000000000000_0001001001001100_1001010100000000"; -- 0.07148104906082153
	pesos_i(1754) := b"1111111111111111_1111111111111111_1110100011010100_1111010001100000"; -- -0.09050057083368301
	pesos_i(1755) := b"0000000000000000_0000000000000000_0001011000011011_0110101000000000"; -- 0.08635580539703369
	pesos_i(1756) := b"1111111111111111_1111111111111111_1100110111101011_1011000110000000"; -- -0.19562235474586487
	pesos_i(1757) := b"0000000000000000_0000000000000000_0010111011111000_0111011001000000"; -- 0.1834787279367447
	pesos_i(1758) := b"0000000000000000_0000000000000000_0001001011001000_1101100001100000"; -- 0.07337715476751328
	pesos_i(1759) := b"1111111111111111_1111111111111111_1101110101001011_1011000001000000"; -- -0.13556383550167084
	pesos_i(1760) := b"0000000000000000_0000000000000000_0000101010010010_1110010110000000"; -- 0.04130396246910095
	pesos_i(1761) := b"1111111111111111_1111111111111111_1111110110000100_0101110111011100"; -- -0.009698995389044285
	pesos_i(1762) := b"0000000000000000_0000000000000000_0101001100101101_1100110100000000"; -- 0.32491761445999146
	pesos_i(1763) := b"0000000000000000_0000000000000000_0010010011000110_1010001111000000"; -- 0.14365600049495697
	pesos_i(1764) := b"1111111111111111_1111111111111111_1110010110111111_0000111000000000"; -- -0.10255348682403564
	pesos_i(1765) := b"0000000000000000_0000000000000000_0101001101101100_1000101100000000"; -- 0.3258749842643738
	pesos_i(1766) := b"0000000000000000_0000000000000000_0001101111001000_0111011011000000"; -- 0.10852758586406708
	pesos_i(1767) := b"0000000000000000_0000000000000000_0111000010010101_1110011000000000"; -- 0.43978726863861084
	pesos_i(1768) := b"0000000000000000_0000000000000000_0011010011001110_1110001101000000"; -- 0.2062818557024002
	pesos_i(1769) := b"0000000000000000_0000000000000000_0010001000100001_0000010010000000"; -- 0.133316308259964
	pesos_i(1770) := b"0000000000000000_0000000000000000_0100101111111100_0111011110000000"; -- 0.29682108759880066
	pesos_i(1771) := b"0000000000000000_0000000000000000_0010000001011101_0001010001000000"; -- 0.1264202743768692
	pesos_i(1772) := b"0000000000000000_0000000000000000_0100110100010001_1101001000000000"; -- 0.30105316638946533
	pesos_i(1773) := b"0000000000000000_0000000000000000_0011101100011000_1100011101000000"; -- 0.2308468371629715
	pesos_i(1774) := b"0000000000000000_0000000000000000_0010101000000101_0011111111000000"; -- 0.16414259374141693
	pesos_i(1775) := b"1111111111111111_1111111111111111_1101111000011111_1100010100000000"; -- -0.13232773542404175
	pesos_i(1776) := b"0000000000000000_0000000000000000_0001110101001111_0100100110000000"; -- 0.11449107527732849
	pesos_i(1777) := b"1111111111111111_1111111111111111_1010100010011011_0110101000000000"; -- -0.3413785696029663
	pesos_i(1778) := b"0000000000000000_0000000000000000_0001001111000111_1111110010100000"; -- 0.07727030664682388
	pesos_i(1779) := b"1111111111111111_1111111111111111_1110111100101101_0100001111100000"; -- -0.06571555882692337
	pesos_i(1780) := b"1111111111111111_1111111111111111_1110110111010110_0101100000000000"; -- -0.07094812393188477
	pesos_i(1781) := b"0000000000000000_0000000000000000_0001001010000000_0010001101100000"; -- 0.07226773351430893
	pesos_i(1782) := b"0000000000000000_0000000000000000_0010010000000111_1101100111000000"; -- 0.14074479043483734
	pesos_i(1783) := b"1111111111111111_1111111111111111_1110010001011110_0000011100000000"; -- -0.10794025659561157
	pesos_i(1784) := b"0000000000000000_0000000000000000_0000110001011011_1100100111000000"; -- 0.048275575041770935
	pesos_i(1785) := b"0000000000000000_0000000000000000_0000000000100010_1001110111010010"; -- 0.0005282056517899036
	pesos_i(1786) := b"0000000000000000_0000000000000000_0000101110100001_1110101000110000"; -- 0.04543937370181084
	pesos_i(1787) := b"1111111111111111_1111111111111111_1111010111100011_1100100011000000"; -- -0.03949303925037384
	pesos_i(1788) := b"0000000000000000_0000000000000000_0000000010010101_0100011001010110"; -- 0.0022777519188821316
	pesos_i(1789) := b"0000000000000000_0000000000000000_0001010110110011_0100101111100000"; -- 0.08476709574460983
	pesos_i(1790) := b"1111111111111111_1111111111111111_1111010001101111_1101110001000000"; -- -0.04516814649105072
	pesos_i(1791) := b"1111111111111111_1111111111111111_1111110111011110_0001100000010100"; -- -0.008329863660037518
	pesos_i(1792) := b"0000000000000000_0000000000000000_0100011000101000_1000100110000000"; -- 0.2740560472011566
	pesos_i(1793) := b"1111111111111111_1111111111111111_1111011000010001_1011011110000000"; -- -0.038792163133621216
	pesos_i(1794) := b"1111111111111111_1111111111111111_1100100010111001_0011010100000000"; -- -0.2159239649772644
	pesos_i(1795) := b"0000000000000000_0000000000000000_0100101001011011_1011101010000000"; -- 0.2904621660709381
	pesos_i(1796) := b"0000000000000000_0000000000000000_0001000011110100_1001100001100000"; -- 0.06623222678899765
	pesos_i(1797) := b"1111111111111111_1111111111111111_0111010100010100_1000110100000000"; -- -0.5426551699638367
	pesos_i(1798) := b"0000000000000000_0000000000000000_0000000110000111_1100001111100010"; -- 0.005977862048894167
	pesos_i(1799) := b"1111111111111111_1111111111111111_1111000000000100_1001000111110000"; -- -0.06243026629090309
	pesos_i(1800) := b"0000000000000000_0000000000000000_0010100011001011_0101101100000000"; -- 0.15935295820236206
	pesos_i(1801) := b"0000000000000000_0000000000000000_0001100111000110_0111010100100000"; -- 0.10068447142839432
	pesos_i(1802) := b"0000000000000000_0000000000000000_0001011010111110_1010000000000000"; -- 0.08884620666503906
	pesos_i(1803) := b"1111111111111111_1111111111111111_1001111001111001_0100011110000000"; -- -0.38096192479133606
	pesos_i(1804) := b"1111111111111111_1111111111111111_1110011011000001_0100000101000000"; -- -0.0986136645078659
	pesos_i(1805) := b"0000000000000000_0000000000000000_0010010110101000_1110000111000000"; -- 0.14710818231105804
	pesos_i(1806) := b"1111111111111111_1111111111111111_1110000111111001_1010111010000000"; -- -0.1172839105129242
	pesos_i(1807) := b"1111111111111111_1111111111111111_1101111100110000_1111010111000000"; -- -0.12815918028354645
	pesos_i(1808) := b"1111111111111111_1111111111111111_1111110000000011_1111000010000100"; -- -0.015564887784421444
	pesos_i(1809) := b"0000000000000000_0000000000000000_0011100100111011_1011100011000000"; -- 0.22356753051280975
	pesos_i(1810) := b"1111111111111111_1111111111111111_1111001010000011_1110011011100000"; -- -0.05267483741044998
	pesos_i(1811) := b"1111111111111111_1111111111111111_1111010010101100_1010111010100000"; -- -0.0442400798201561
	pesos_i(1812) := b"0000000000000000_0000000000000000_0001000110010001_1001100001100000"; -- 0.06862785667181015
	pesos_i(1813) := b"0000000000000000_0000000000000000_0001010011010101_1011011011000000"; -- 0.0813860148191452
	pesos_i(1814) := b"1111111111111111_1111111111111111_1110010000100101_1100010011000000"; -- -0.10879869759082794
	pesos_i(1815) := b"1111111111111111_1111111111111111_1100011111011100_0111101100000000"; -- -0.21929198503494263
	pesos_i(1816) := b"1111111111111111_1111111111111111_1110110110111011_1111010111100000"; -- -0.07135070115327835
	pesos_i(1817) := b"1111111111111111_1111111111111111_1111101110001011_1101011011101000"; -- -0.01739746890962124
	pesos_i(1818) := b"1111111111111111_1111111111111111_1101001110111111_0100101110000000"; -- -0.17286232113838196
	pesos_i(1819) := b"0000000000000000_0000000000000000_0011001000101111_1100101000000000"; -- 0.19604170322418213
	pesos_i(1820) := b"1111111111111111_1111111111111111_1100000101110110_1101011000000000"; -- -0.24428045749664307
	pesos_i(1821) := b"0000000000000000_0000000000000000_0011001110001101_1101100000000000"; -- 0.20138311386108398
	pesos_i(1822) := b"1111111111111111_1111111111111111_1101010010101011_1001001011000000"; -- -0.1692570000886917
	pesos_i(1823) := b"1111111111111111_1111111111111111_1101000000011100_0101111001000000"; -- -0.18706713616847992
	pesos_i(1824) := b"0000000000000000_0000000000000000_0010011111100011_1110001101000000"; -- 0.1558210402727127
	pesos_i(1825) := b"0000000000000000_0000000000000000_0010110100001100_1011101010000000"; -- 0.1759754717350006
	pesos_i(1826) := b"0000000000000000_0000000000000000_0000000010101000_1000101000000100"; -- 0.0025717029348015785
	pesos_i(1827) := b"0000000000000000_0000000000000000_0001100000101010_1001101100100000"; -- 0.09440011531114578
	pesos_i(1828) := b"0000000000000000_0000000000000000_0010111101000100_0000111100000000"; -- 0.18463224172592163
	pesos_i(1829) := b"0000000000000000_0000000000000000_0010001100110110_1101111000000000"; -- 0.13755595684051514
	pesos_i(1830) := b"1111111111111111_1111111111111111_1110101111101001_0111101101100000"; -- -0.07846859842538834
	pesos_i(1831) := b"0000000000000000_0000000000000000_0001010111000100_1011101000000000"; -- 0.08503305912017822
	pesos_i(1832) := b"0000000000000000_0000000000000000_0101111110000110_0000001010000000"; -- 0.37313857674598694
	pesos_i(1833) := b"1111111111111111_1111111111111111_1110111101011101_1010001111100000"; -- -0.06497741490602493
	pesos_i(1834) := b"1111111111111111_1111111111111111_1100100111010001_1011111001000000"; -- -0.21164332330226898
	pesos_i(1835) := b"1111111111111111_1111111111111111_1001001001011111_0001110100000000"; -- -0.428236186504364
	pesos_i(1836) := b"1111111111111111_1111111111111111_1010110101101000_0100110000000000"; -- -0.32262730598449707
	pesos_i(1837) := b"0000000000000000_0000000000000000_0001011011000001_1011010100100000"; -- 0.08889324218034744
	pesos_i(1838) := b"1111111111111111_1111111111111111_1111101011000011_0010101110001000"; -- -0.02045944146811962
	pesos_i(1839) := b"0000000000000000_0000000000000000_0100110100101000_0111001000000000"; -- 0.3013983964920044
	pesos_i(1840) := b"0000000000000000_0000000000000000_0010000110111111_1110101111000000"; -- 0.1318347305059433
	pesos_i(1841) := b"1111111111111111_1111111111111111_1100111110111011_1101011000000000"; -- -0.18854010105133057
	pesos_i(1842) := b"0000000000000000_0000000000000000_0001000100001001_1001010111100000"; -- 0.06655251234769821
	pesos_i(1843) := b"0000000000000000_0000000000000000_0000111011110000_1110000111000000"; -- 0.058363065123558044
	pesos_i(1844) := b"0000000000000000_0000000000000000_0001111011100011_1100111011100000"; -- 0.12066357582807541
	pesos_i(1845) := b"1111111111111111_1111111111111111_1110000010010111_1011111000000000"; -- -0.12268459796905518
	pesos_i(1846) := b"0000000000000000_0000000000000000_0011000000111010_0010100011000000"; -- 0.1883874386548996
	pesos_i(1847) := b"1111111111111111_1111111111111111_1110101011010010_0001111110100000"; -- -0.08273126929998398
	pesos_i(1848) := b"0000000000000000_0000000000000000_0100110010101000_0110011010000000"; -- 0.2994445860385895
	pesos_i(1849) := b"0000000000000000_0000000000000000_0000011011100011_1100011110110000"; -- 0.026913147419691086
	pesos_i(1850) := b"1111111111111111_1111111111111111_1111100010111111_0000001000000000"; -- -0.02833545207977295
	pesos_i(1851) := b"0000000000000000_0000000000000000_0001011000011011_1101011001100000"; -- 0.08636226505041122
	pesos_i(1852) := b"1111111111111111_1111111111111111_1101011110010010_0111001110000000"; -- -0.15792158246040344
	pesos_i(1853) := b"0000000000000000_0000000000000000_0010000010000010_0011010101000000"; -- 0.1269868165254593
	pesos_i(1854) := b"0000000000000000_0000000000000000_0001100100010010_0101001010100000"; -- 0.09793583303689957
	pesos_i(1855) := b"1111111111111111_1111111111111111_1101111100111100_1110100000000000"; -- -0.1279768943786621
	pesos_i(1856) := b"0000000000000000_0000000000000000_0010110100111010_0000101100000000"; -- 0.17666691541671753
	pesos_i(1857) := b"0000000000000000_0000000000000000_0010101010100000_1000110010000000"; -- 0.16651228070259094
	pesos_i(1858) := b"0000000000000000_0000000000000000_0011010000000011_0001111100000000"; -- 0.20317262411117554
	pesos_i(1859) := b"0000000000000000_0000000000000000_0000010110010000_1010100010110000"; -- 0.02173857018351555
	pesos_i(1860) := b"0000000000000000_0000000000000000_0000110011001011_1111100011110000"; -- 0.049987372010946274
	pesos_i(1861) := b"0000000000000000_0000000000000000_0000001010100101_0100010010011100"; -- 0.010334289632737637
	pesos_i(1862) := b"1111111111111111_1111111111111111_1110111001101000_0111001000100000"; -- -0.06871878355741501
	pesos_i(1863) := b"0000000000000000_0000000000000000_0000000011110100_0000011010011011"; -- 0.0037235382478684187
	pesos_i(1864) := b"0000000000000000_0000000000000000_0001110101110100_1111110010100000"; -- 0.11506632715463638
	pesos_i(1865) := b"0000000000000000_0000000000000000_0001111101000010_0010100010000000"; -- 0.1221032440662384
	pesos_i(1866) := b"1111111111111111_1111111111111111_1111110101101100_1111001100001000"; -- -0.01005631498992443
	pesos_i(1867) := b"1111111111111111_1111111111111111_1110110001111010_1101111010100000"; -- -0.07625015825033188
	pesos_i(1868) := b"1111111111111111_1111111111111111_1111000100000011_1001111001100000"; -- -0.0585385337471962
	pesos_i(1869) := b"1111111111111111_1111111111111111_1101101111010100_0001100010000000"; -- -0.141294926404953
	pesos_i(1870) := b"1111111111111111_1111111111111111_1110111100001101_0010101101100000"; -- -0.06620530039072037
	pesos_i(1871) := b"0000000000000000_0000000000000000_0000011001000001_1000111111010000"; -- 0.02443789318203926
	pesos_i(1872) := b"1111111111111111_1111111111111111_1101111011010101_1100101011000000"; -- -0.1295502930879593
	pesos_i(1873) := b"0000000000000000_0000000000000000_0001100010110010_0000100011000000"; -- 0.09646658599376678
	pesos_i(1874) := b"0000000000000000_0000000000000000_0100000011010000_0011010110000000"; -- 0.2531770169734955
	pesos_i(1875) := b"0000000000000000_0000000000000000_0010101000101111_0101011111000000"; -- 0.16478489339351654
	pesos_i(1876) := b"0000000000000000_0000000000000000_0010111011010110_1101000101000000"; -- 0.18296535313129425
	pesos_i(1877) := b"0000000000000000_0000000000000000_0010101010011100_0110000100000000"; -- 0.1664486527442932
	pesos_i(1878) := b"1111111111111111_1111111111111111_1111111101101101_1011000001101110"; -- -0.0022325259633362293
	pesos_i(1879) := b"1111111111111111_1111111111111111_1111000011101001_0011111011000000"; -- -0.058940961956977844
	pesos_i(1880) := b"1111111111111111_1111111111111111_1111010000011110_1011101011110000"; -- -0.0464060939848423
	pesos_i(1881) := b"0000000000000000_0000000000000000_0000100110111001_1100001000110000"; -- 0.03799070045351982
	pesos_i(1882) := b"0000000000000000_0000000000000000_0000011011100011_0011011100111000"; -- 0.02690453641116619
	pesos_i(1883) := b"1111111111111111_1111111111111111_1111010000111000_0101100001010000"; -- -0.04601524397730827
	pesos_i(1884) := b"1111111111111111_1111111111111111_1110101001010000_1010010011100000"; -- -0.08470696955919266
	pesos_i(1885) := b"0000000000000000_0000000000000000_0000001010101010_1110101001010100"; -- 0.010420461185276508
	pesos_i(1886) := b"1111111111111111_1111111111111111_1101111001011110_1110010111000000"; -- -0.13136447966098785
	pesos_i(1887) := b"1111111111111111_1111111111111111_1101111001111111_1110100111000000"; -- -0.13086070120334625
	pesos_i(1888) := b"1111111111111111_1111111111111111_1110011101010001_0101000110100000"; -- -0.09641542285680771
	pesos_i(1889) := b"1111111111111111_1111111111111111_1110100111011001_0010001101000000"; -- -0.08653049170970917
	pesos_i(1890) := b"1111111111111111_1111111111111111_1110011001101100_1001110000100000"; -- -0.09990524500608444
	pesos_i(1891) := b"1111111111111111_1111111111111111_1111011111100000_0111001001000000"; -- -0.03173147141933441
	pesos_i(1892) := b"1111111111111111_1111111111111111_1001110101101110_0001111100000000"; -- -0.38503843545913696
	pesos_i(1893) := b"0000000000000000_0000000000000000_0000011000001110_1100111111001000"; -- 0.023663507774472237
	pesos_i(1894) := b"0000000000000000_0000000000000000_0011111001110001_0010000101000000"; -- 0.24391372501850128
	pesos_i(1895) := b"0000000000000000_0000000000000000_0001110011010010_1000110100000000"; -- 0.11258774995803833
	pesos_i(1896) := b"1111111111111111_1111111111111111_1101111100000011_0100011010000000"; -- -0.12885627150535583
	pesos_i(1897) := b"0000000000000000_0000000000000000_0011010010001100_1101011110000000"; -- 0.2052740752696991
	pesos_i(1898) := b"0000000000000000_0000000000000000_0010001011101101_0101000111000000"; -- 0.1364337056875229
	pesos_i(1899) := b"0000000000000000_0000000000000000_0000111001011010_0010101110110000"; -- 0.056063394993543625
	pesos_i(1900) := b"0000000000000000_0000000000000000_0011101000011101_1110111011000000"; -- 0.22701923549175262
	pesos_i(1901) := b"0000000000000000_0000000000000000_0001011000011010_0101010000000000"; -- 0.08633923530578613
	pesos_i(1902) := b"0000000000000000_0000000000000000_0000111111001101_1110011010000000"; -- 0.06173554062843323
	pesos_i(1903) := b"0000000000000000_0000000000000000_0000100011010000_0101100111010000"; -- 0.03442918136715889
	pesos_i(1904) := b"0000000000000000_0000000000000000_0010100001111111_1101011111000000"; -- 0.1582007259130478
	pesos_i(1905) := b"1111111111111111_1111111111111111_1100110000100101_1110100110000000"; -- -0.20254650712013245
	pesos_i(1906) := b"1111111111111111_1111111111111111_1110101010000011_0001100001000000"; -- -0.0839371532201767
	pesos_i(1907) := b"0000000000000000_0000000000000000_0000110011010111_0110001001010000"; -- 0.05016149953007698
	pesos_i(1908) := b"0000000000000000_0000000000000000_0010111011101111_0011011001000000"; -- 0.18333758413791656
	pesos_i(1909) := b"0000000000000000_0000000000000000_0001010001010001_1111011010000000"; -- 0.07937565445899963
	pesos_i(1910) := b"1111111111111111_1111111111111111_1111001100111100_0110001111000000"; -- -0.049859777092933655
	pesos_i(1911) := b"1111111111111111_1111111111111111_1101010000100100_1111110001000000"; -- -0.1713106483221054
	pesos_i(1912) := b"1111111111111111_1111111111111111_1111001011001000_1100010011110000"; -- -0.051624003797769547
	pesos_i(1913) := b"0000000000000000_0000000000000000_0000011111010011_0101100011001000"; -- 0.030568646267056465
	pesos_i(1914) := b"0000000000000000_0000000000000000_0000110001011011_1100101111010000"; -- 0.048275697976350784
	pesos_i(1915) := b"1111111111111111_1111111111111111_1111110000001111_1111111010000000"; -- -0.015380948781967163
	pesos_i(1916) := b"0000000000000000_0000000000000000_0000101011100110_1101101000110000"; -- 0.04258502647280693
	pesos_i(1917) := b"1111111111111111_1111111111111111_1010100010000101_1011110110000000"; -- -0.34170928597450256
	pesos_i(1918) := b"1111111111111111_1111111111111111_1100110101010000_0010000111000000"; -- -0.19799603521823883
	pesos_i(1919) := b"0000000000000000_0000000000000000_0000001000100000_1000101011011000"; -- 0.008309056982398033
	pesos_i(1920) := b"1111111111111111_1111111111111111_1111101110111001_0001100001000000"; -- -0.016706928610801697
	pesos_i(1921) := b"1111111111111111_1111111111111111_1110011010001011_0010000011100000"; -- -0.09943956881761551
	pesos_i(1922) := b"1111111111111111_1111111111111111_1100110110110101_0011010000000000"; -- -0.19645380973815918
	pesos_i(1923) := b"0000000000000000_0000000000000000_0010101110101111_0110110111000000"; -- 0.1706455796957016
	pesos_i(1924) := b"0000000000000000_0000000000000000_0000010101101000_1000110101110000"; -- 0.02112659439444542
	pesos_i(1925) := b"1111111111111111_1111111111111111_1011001011001110_1101011010000000"; -- -0.3015314042568207
	pesos_i(1926) := b"1111111111111111_1111111111111111_1111111110100101_1100101110001110"; -- -0.001376416883431375
	pesos_i(1927) := b"1111111111111111_1111111111111111_1111000010111011_1100001011010000"; -- -0.059634994715452194
	pesos_i(1928) := b"0000000000000000_0000000000000000_0001001101101010_1001011010100000"; -- 0.0758451595902443
	pesos_i(1929) := b"0000000000000000_0000000000000000_0010010000101011_0011111111000000"; -- 0.14128492772579193
	pesos_i(1930) := b"0000000000000000_0000000000000000_0010000010110000_1001001010000000"; -- 0.1276942789554596
	pesos_i(1931) := b"1111111111111111_1111111111111111_1011101100101011_1110100110000000"; -- -0.26886120438575745
	pesos_i(1932) := b"0000000000000000_0000000000000000_0010001101001110_1101000100000000"; -- 0.13792139291763306
	pesos_i(1933) := b"0000000000000000_0000000000000000_0000001011001011_0011111011010000"; -- 0.010913778096437454
	pesos_i(1934) := b"1111111111111111_1111111111111111_1101111111010100_1010011001000000"; -- -0.1256614774465561
	pesos_i(1935) := b"1111111111111111_1111111111111111_1110010111010101_0111101010000000"; -- -0.10221132636070251
	pesos_i(1936) := b"1111111111111111_1111111111111111_1110100101101011_1101101000000000"; -- -0.08819806575775146
	pesos_i(1937) := b"0000000000000000_0000000000000000_0010101110111011_1101100010000000"; -- 0.17083504796028137
	pesos_i(1938) := b"1111111111111111_1111111111111111_1100111111011000_0111011100000000"; -- -0.18810325860977173
	pesos_i(1939) := b"1111111111111111_1111111111111111_1110010100001001_0011100110100000"; -- -0.10532798618078232
	pesos_i(1940) := b"0000000000000000_0000000000000000_0010111000100000_0111000011000000"; -- 0.18018250167369843
	pesos_i(1941) := b"0000000000000000_0000000000000000_0000001011100110_1111011100000000"; -- 0.011336743831634521
	pesos_i(1942) := b"1111111111111111_1111111111111111_1110000010010000_0100100010100000"; -- -0.12279840558767319
	pesos_i(1943) := b"0000000000000000_0000000000000000_0001101000011011_0111010111100000"; -- 0.1019815132021904
	pesos_i(1944) := b"1111111111111111_1111111111111111_1101000000101011_0001111001000000"; -- -0.18684206902980804
	pesos_i(1945) := b"0000000000000000_0000000000000000_0010100010011111_0111101011000000"; -- 0.15868346393108368
	pesos_i(1946) := b"1111111111111111_1111111111111111_1011001011110110_0000001110000000"; -- -0.3009336292743683
	pesos_i(1947) := b"1111111111111111_1111111111111111_1110010101010110_1111001101000000"; -- -0.10414199531078339
	pesos_i(1948) := b"1111111111111111_1111111111111111_0110000010100110_1101110100000000"; -- -0.6224538683891296
	pesos_i(1949) := b"0000000000000000_0000000000000000_0010111010001111_0000001010000000"; -- 0.18186965584754944
	pesos_i(1950) := b"1111111111111111_1111111111111111_1101011101010111_0100111110000000"; -- -0.15882399678230286
	pesos_i(1951) := b"1111111111111111_1111111111111111_1110000111111111_0101110011000000"; -- -0.11719723045825958
	pesos_i(1952) := b"0000000000000000_0000000000000000_0010101011000010_1101111110000000"; -- 0.1670360267162323
	pesos_i(1953) := b"0000000000000000_0000000000000000_0000001100100000_0101010001010100"; -- 0.0122120575979352
	pesos_i(1954) := b"1111111111111111_1111111111111111_1110001010111111_0100011111100000"; -- -0.11426878720521927
	pesos_i(1955) := b"1111111111111111_1111111111111111_1111011101010100_1111111101000000"; -- -0.03385929763317108
	pesos_i(1956) := b"0000000000000000_0000000000000000_0011000110000111_0101101100000000"; -- 0.19347161054611206
	pesos_i(1957) := b"0000000000000000_0000000000000000_0100111100001111_1011001010000000"; -- 0.3088332712650299
	pesos_i(1958) := b"0000000000000000_0000000000000000_0000101100110000_0101111010010000"; -- 0.04370680823922157
	pesos_i(1959) := b"1111111111111111_1111111111111111_1110101001000011_0100000100000000"; -- -0.0849112868309021
	pesos_i(1960) := b"0000000000000000_0000000000000000_0011011101101110_1001101101000000"; -- 0.21653147041797638
	pesos_i(1961) := b"1111111111111111_1111111111111111_1110001100001010_1100011110100000"; -- -0.11311676353216171
	pesos_i(1962) := b"1111111111111111_1111111111111111_1101101100111100_1011111111000000"; -- -0.14360429346561432
	pesos_i(1963) := b"1111111111111111_1111111111111111_1011110000010001_1010011100000000"; -- -0.26535564661026
	pesos_i(1964) := b"1111111111111111_1111111111111111_1110011100011000_0110110001000000"; -- -0.09728358685970306
	pesos_i(1965) := b"0000000000000000_0000000000000000_0000100100001000_0101000000000000"; -- 0.03528308868408203
	pesos_i(1966) := b"1111111111111111_1111111111111111_1110000011101010_0110001001100000"; -- -0.12142357975244522
	pesos_i(1967) := b"0000000000000000_0000000000000000_0000100100100011_1010011111100000"; -- 0.03570031374692917
	pesos_i(1968) := b"0000000000000000_0000000000000000_0000000110110000_1010101111101010"; -- 0.006602043751627207
	pesos_i(1969) := b"1111111111111111_1111111111111111_1010110100000110_0011100000000000"; -- -0.3241238594055176
	pesos_i(1970) := b"1111111111111111_1111111111111111_1111000101111001_1011111100000000"; -- -0.0567360520362854
	pesos_i(1971) := b"1111111111111111_1111111111111111_1111001001110100_1010001000000000"; -- -0.05290782451629639
	pesos_i(1972) := b"1111111111111111_1111111111111111_1111001000000011_1001110100100000"; -- -0.05463235825300217
	pesos_i(1973) := b"0000000000000000_0000000000000000_0001101000001000_1111110100100000"; -- 0.10169965773820877
	pesos_i(1974) := b"0000000000000000_0000000000000000_0100001010011001_1011011000000000"; -- 0.2601579427719116
	pesos_i(1975) := b"1111111111111111_1111111111111111_1001011101101001_1101110010000000"; -- -0.4085409343242645
	pesos_i(1976) := b"0000000000000000_0000000000000000_0000111000011110_0000010011110000"; -- 0.05514555796980858
	pesos_i(1977) := b"0000000000000000_0000000000000000_0000000011110111_0111111100100110"; -- 0.0037764995358884335
	pesos_i(1978) := b"1111111111111111_1111111111111111_1111001001110000_1101010010000000"; -- -0.05296584963798523
	pesos_i(1979) := b"1111111111111111_1111111111111111_1111111101001100_1010011000001110"; -- -0.002736684400588274
	pesos_i(1980) := b"1111111111111111_1111111111111111_1011110001101001_0001101000000000"; -- -0.26402127742767334
	pesos_i(1981) := b"0000000000000000_0000000000000000_0001001111001100_0001001111000000"; -- 0.07733272016048431
	pesos_i(1982) := b"1111111111111111_1111111111111111_1101001000110001_1100100011000000"; -- -0.17892785370349884
	pesos_i(1983) := b"1111111111111111_1111111111111111_0111100010000110_1000110100000000"; -- -0.5291969180107117
	pesos_i(1984) := b"0000000000000000_0000000000000000_0011000111001011_0100010000000000"; -- 0.19450783729553223
	pesos_i(1985) := b"0000000000000000_0000000000000000_0001111110100110_0001110011000000"; -- 0.12362842261791229
	pesos_i(1986) := b"0000000000000000_0000000000000000_0001011101111000_1000111001100000"; -- 0.0916832908987999
	pesos_i(1987) := b"0000000000000000_0000000000000000_0001000111011100_0100101010000000"; -- 0.06976762413978577
	pesos_i(1988) := b"1111111111111111_1111111111111111_1010100101101011_0100000000000000"; -- -0.3382072448730469
	pesos_i(1989) := b"1111111111111111_1111111111111111_1101111010110011_1100000001000000"; -- -0.13006971776485443
	pesos_i(1990) := b"0000000000000000_0000000000000000_0011100000000011_1000011101000000"; -- 0.21880383789539337
	pesos_i(1991) := b"0000000000000000_0000000000000000_0001011010010011_0001011011000000"; -- 0.08818189799785614
	pesos_i(1992) := b"1111111111111111_1111111111111111_1111011101100110_0100110000010000"; -- -0.03359531983733177
	pesos_i(1993) := b"0000000000000000_0000000000000000_0000011011011000_1010101010010000"; -- 0.026743564754724503
	pesos_i(1994) := b"1111111111111111_1111111111111111_1110100111001110_0001011001100000"; -- -0.08669910579919815
	pesos_i(1995) := b"0000000000000000_0000000000000000_0001100000110000_1010001111000000"; -- 0.09449218213558197
	pesos_i(1996) := b"1111111111111111_1111111111111111_1110010101011111_0011100101100000"; -- -0.10401574522256851
	pesos_i(1997) := b"1111111111111111_1111111111111111_1100111011000100_1110011110000000"; -- -0.1923079788684845
	pesos_i(1998) := b"0000000000000000_0000000000000000_0010000000110101_1111001010000000"; -- 0.12582316994667053
	pesos_i(1999) := b"1111111111111111_1111111111111111_1011010101101101_0110111010000000"; -- -0.2912989556789398
	pesos_i(2000) := b"1111111111111111_1111111111111111_1110001110001110_1001000110100000"; -- -0.11110582202672958
	pesos_i(2001) := b"0000000000000000_0000000000000000_0010000110110011_0100101100000000"; -- 0.13164204359054565
	pesos_i(2002) := b"0000000000000000_0000000000000000_0000110001011100_1000101000000000"; -- 0.048287034034729004
	pesos_i(2003) := b"0000000000000000_0000000000000000_0011011011100001_1111000011000000"; -- 0.21438507735729218
	pesos_i(2004) := b"0000000000000000_0000000000000000_0000101010110000_0011001010000000"; -- 0.04175105690956116
	pesos_i(2005) := b"0000000000000000_0000000000000000_0000001000011110_1110001100001100"; -- 0.008283796720206738
	pesos_i(2006) := b"1111111111111111_1111111111111111_1111110000010110_0101100011100100"; -- -0.015284008346498013
	pesos_i(2007) := b"1111111111111111_1111111111111111_1100111000110101_0011011001000000"; -- -0.19450055062770844
	pesos_i(2008) := b"1111111111111111_1111111111111111_1110000101100001_1001111010000000"; -- -0.1196042001247406
	pesos_i(2009) := b"0000000000000000_0000000000000000_0011101110110011_1010001110000000"; -- 0.23320981860160828
	pesos_i(2010) := b"0000000000000000_0000000000000000_0000001100101111_0010010110011000"; -- 0.012438153848052025
	pesos_i(2011) := b"0000000000000000_0000000000000000_0000101100110010_1010110010010000"; -- 0.04374197497963905
	pesos_i(2012) := b"0000000000000000_0000000000000000_0000110000010000_1101100010110000"; -- 0.04713205620646477
	pesos_i(2013) := b"1111111111111111_1111111111111111_1101100111011110_1011000111000000"; -- -0.14894570410251617
	pesos_i(2014) := b"1111111111111111_1111111111111111_1111001011110000_1010010111100000"; -- -0.05101550370454788
	pesos_i(2015) := b"1111111111111111_1111111111111111_1100101110010001_1101011010000000"; -- -0.20480594038963318
	pesos_i(2016) := b"0000000000000000_0000000000000000_0001111110111101_0111010001000000"; -- 0.12398459017276764
	pesos_i(2017) := b"1111111111111111_1111111111111111_1101011000110001_0110100111000000"; -- -0.1633085161447525
	pesos_i(2018) := b"1111111111111111_1111111111111111_1100000011100101_1111001111000000"; -- -0.2464912086725235
	pesos_i(2019) := b"0000000000000000_0000000000000000_0010110000110111_1001010010000000"; -- 0.17272308468818665
	pesos_i(2020) := b"1111111111111111_1111111111111111_1000111011001010_0001001000000000"; -- -0.44222915172576904
	pesos_i(2021) := b"1111111111111111_1111111111111111_1101101100110101_1100000000000000"; -- -0.14371109008789062
	pesos_i(2022) := b"0000000000000000_0000000000000000_0101100111000001_0111000100000000"; -- 0.3506079316139221
	pesos_i(2023) := b"1111111111111111_1111111111111111_1111100100101111_1000010110001000"; -- -0.026618627831339836
	pesos_i(2024) := b"0000000000000000_0000000000000000_0011001010100011_1000110011000000"; -- 0.19780807197093964
	pesos_i(2025) := b"0000000000000000_0000000000000000_0001100110110010_1010011010000000"; -- 0.1003822386264801
	pesos_i(2026) := b"0000000000000000_0000000000000000_0010010001011011_0110000111000000"; -- 0.1420193761587143
	pesos_i(2027) := b"1111111111111111_1111111111111111_1110011001001010_0101100100100000"; -- -0.1004280373454094
	pesos_i(2028) := b"0000000000000000_0000000000000000_0001001110010110_1000000001000000"; -- 0.07651521265506744
	pesos_i(2029) := b"0000000000000000_0000000000000000_0000100011010001_0110001101010000"; -- 0.034445006400346756
	pesos_i(2030) := b"1111111111111111_1111111111111111_1100011100000110_1001101001000000"; -- -0.2225555032491684
	pesos_i(2031) := b"1111111111111111_1111111111111111_1111101010010000_0001110110011000"; -- -0.02123847045004368
	pesos_i(2032) := b"0000000000000000_0000000000000000_0011000110001011_1110000100000000"; -- 0.19354063272476196
	pesos_i(2033) := b"1111111111111111_1111111111111111_1011100111011111_0101011110000000"; -- -0.27393582463264465
	pesos_i(2034) := b"0000000000000000_0000000000000000_0001111110010110_0000100110000000"; -- 0.12338313460350037
	pesos_i(2035) := b"1111111111111111_1111111111111111_1110011101001001_0011110110100000"; -- -0.09653868526220322
	pesos_i(2036) := b"0000000000000000_0000000000000000_0100110011001000_1001001010000000"; -- 0.2999354898929596
	pesos_i(2037) := b"1111111111111111_1111111111111111_1110010011100100_0110100101100000"; -- -0.1058897152543068
	pesos_i(2038) := b"1111111111111111_1111111111111111_1110111101010000_0010100011000000"; -- -0.0651831179857254
	pesos_i(2039) := b"1111111111111111_1111111111111111_1110110010110001_1001101100100000"; -- -0.07541494816541672
	pesos_i(2040) := b"0000000000000000_0000000000000000_0001101000100000_0110010111100000"; -- 0.10205685347318649
	pesos_i(2041) := b"1111111111111111_1111111111111111_1110000010001010_1100000000100000"; -- -0.12288283556699753
	pesos_i(2042) := b"0000000000000000_0000000000000000_0010011010011101_1111101100000000"; -- 0.15084809064865112
	pesos_i(2043) := b"1111111111111111_1111111111111111_1110000100101110_0100101110000000"; -- -0.12038734555244446
	pesos_i(2044) := b"1111111111111111_1111111111111111_1110100110110100_0011011110100000"; -- -0.08709385246038437
	pesos_i(2045) := b"0000000000000000_0000000000000000_0001010011001110_1010001011000000"; -- 0.0812780112028122
	pesos_i(2046) := b"1111111111111111_1111111111111111_1011111001101011_1011010010000000"; -- -0.25616905093193054
	pesos_i(2047) := b"1111111111111111_1111111111111111_1100000110011011_0110101111000000"; -- -0.24372221529483795
	pesos_i(2048) := b"1111111111111111_1111111111111111_1110110001100001_0111110000100000"; -- -0.07663749903440475
	pesos_i(2049) := b"0000000000000000_0000000000000000_0000110111100010_0101100010000000"; -- 0.05423501133918762
	pesos_i(2050) := b"1111111111111111_1111111111111111_1111111110111000_0010010010010100"; -- -0.0010964524699375033
	pesos_i(2051) := b"1111111111111111_1111111111111111_1111111001001010_1101100011100010"; -- -0.00667042238637805
	pesos_i(2052) := b"0000000000000000_0000000000000000_0000100011001101_0100110000000000"; -- 0.03438258171081543
	pesos_i(2053) := b"1111111111111111_1111111111111111_1111100010011110_1111110110100000"; -- -0.02882399410009384
	pesos_i(2054) := b"0000000000000000_0000000000000000_0000100101100010_1001101010110000"; -- 0.03666083142161369
	pesos_i(2055) := b"0000000000000000_0000000000000000_0000101001000101_1001110101000000"; -- 0.04012472927570343
	pesos_i(2056) := b"0000000000000000_0000000000000000_0001001001111000_0011111100100000"; -- 0.07214731723070145
	pesos_i(2057) := b"1111111111111111_1111111111111111_1011001000111000_1111110110000000"; -- -0.30381789803504944
	pesos_i(2058) := b"0000000000000000_0000000000000000_0010011101011000_1111110100000000"; -- 0.15370160341262817
	pesos_i(2059) := b"0000000000000000_0000000000000000_0011000110101111_0111100110000000"; -- 0.1940837800502777
	pesos_i(2060) := b"0000000000000000_0000000000000000_0000100111100110_1110011010110000"; -- 0.03867952153086662
	pesos_i(2061) := b"1111111111111111_1111111111111111_1111011101101100_0010010011100000"; -- -0.03350610285997391
	pesos_i(2062) := b"0000000000000000_0000000000000000_0100110110001100_1011100110000000"; -- 0.30292853713035583
	pesos_i(2063) := b"0000000000000000_0000000000000000_0010100011011001_0110010010000000"; -- 0.15956714749336243
	pesos_i(2064) := b"1111111111111111_1111111111111111_1010010100001110_0110000110000000"; -- -0.3552493155002594
	pesos_i(2065) := b"1111111111111111_1111111111111111_1111001001011111_0000000101110000"; -- -0.053237829357385635
	pesos_i(2066) := b"1111111111111111_1111111111111111_1111111011110110_0000000001101100"; -- -0.004058812744915485
	pesos_i(2067) := b"0000000000000000_0000000000000000_0011101011111010_0111100010000000"; -- 0.23038437962532043
	pesos_i(2068) := b"0000000000000000_0000000000000000_0001100010010001_1111111010100000"; -- 0.09597770124673843
	pesos_i(2069) := b"0000000000000000_0000000000000000_0001101000001100_1010000001000000"; -- 0.10175515711307526
	pesos_i(2070) := b"0000000000000000_0000000000000000_0011000110100011_1011110111000000"; -- 0.19390474259853363
	pesos_i(2071) := b"1111111111111111_1111111111111111_1011110111101101_0010100000000000"; -- -0.2581000328063965
	pesos_i(2072) := b"0000000000000000_0000000000000000_0000000011100001_1001101000010000"; -- 0.0034424103796482086
	pesos_i(2073) := b"0000000000000000_0000000000000000_0000011000110101_1110100010011000"; -- 0.024260079488158226
	pesos_i(2074) := b"0000000000000000_0000000000000000_0001010000101001_1010000101100000"; -- 0.07876022905111313
	pesos_i(2075) := b"1111111111111111_1111111111111111_1011001110010011_0100101000000000"; -- -0.2985337972640991
	pesos_i(2076) := b"0000000000000000_0000000000000000_0010000001110000_0000110110000000"; -- 0.12670978903770447
	pesos_i(2077) := b"1111111111111111_1111111111111111_1111101011111010_0101010000110000"; -- -0.019617784768342972
	pesos_i(2078) := b"1111111111111111_1111111111111111_1111110000000110_0001001001010000"; -- -0.01553235575556755
	pesos_i(2079) := b"1111111111111111_1111111111111111_1111000010101010_0000000011000000"; -- -0.05990596115589142
	pesos_i(2080) := b"0000000000000000_0000000000000000_0100000010000101_1011010010000000"; -- 0.25204017758369446
	pesos_i(2081) := b"1111111111111111_1111111111111111_1101110110100011_0001010001000000"; -- -0.1342303603887558
	pesos_i(2082) := b"1111111111111111_1111111111111111_1111100011101000_1101101001111000"; -- -0.027696939185261726
	pesos_i(2083) := b"0000000000000000_0000000000000000_0000101000110000_0010001000000000"; -- 0.03979694843292236
	pesos_i(2084) := b"1111111111111111_1111111111111111_1111011001000111_0110111100010000"; -- -0.03797250613570213
	pesos_i(2085) := b"0000000000000000_0000000000000000_0000111000000110_1011001010010000"; -- 0.054789695888757706
	pesos_i(2086) := b"1111111111111111_1111111111111111_1010110100100001_0001000010000000"; -- -0.3237142264842987
	pesos_i(2087) := b"1111111111111111_1111111111111111_1111010111100001_0110101100000000"; -- -0.03952914476394653
	pesos_i(2088) := b"1111111111111111_1111111111111111_1110100011111000_0010111111000000"; -- -0.08996297419071198
	pesos_i(2089) := b"0000000000000000_0000000000000000_0000000011111010_0110110110011101"; -- 0.0038212307263165712
	pesos_i(2090) := b"0000000000000000_0000000000000000_0110011100110000_0011010110000000"; -- 0.4030793607234955
	pesos_i(2091) := b"0000000000000000_0000000000000000_0000011101110100_0110011001111000"; -- 0.02911987714469433
	pesos_i(2092) := b"0000000000000000_0000000000000000_0100010000000100_0110100010000000"; -- 0.26569226384162903
	pesos_i(2093) := b"0000000000000000_0000000000000000_0001100001000001_0101100000000000"; -- 0.09474706649780273
	pesos_i(2094) := b"0000000000000000_0000000000000000_0000000111010100_0111011010001000"; -- 0.007148178294301033
	pesos_i(2095) := b"0000000000000000_0000000000000000_0000000101101101_1011110011101100"; -- 0.005580718629062176
	pesos_i(2096) := b"0000000000000000_0000000000000000_0000110111010110_0101011111000000"; -- 0.05405186116695404
	pesos_i(2097) := b"1111111111111111_1111111111111111_1111101011110010_0111011011011000"; -- -0.019737789407372475
	pesos_i(2098) := b"1111111111111111_1111111111111111_1100010100101011_1011100101000000"; -- -0.22980158030986786
	pesos_i(2099) := b"1111111111111111_1111111111111111_1111000001000111_0001010100110000"; -- -0.06141536310315132
	pesos_i(2100) := b"1111111111111111_1111111111111111_1100010011111110_1000001001000000"; -- -0.230491504073143
	pesos_i(2101) := b"1111111111111111_1111111111111111_1111001011000001_0100001111010000"; -- -0.05173851177096367
	pesos_i(2102) := b"1111111111111111_1111111111111111_1101000010110111_1110111000000000"; -- -0.18469345569610596
	pesos_i(2103) := b"0000000000000000_0000000000000000_0001101100111111_1000101010000000"; -- 0.10643830895423889
	pesos_i(2104) := b"1111111111111111_1111111111111111_1101011110001110_0000100010000000"; -- -0.1579889953136444
	pesos_i(2105) := b"0000000000000000_0000000000000000_0100100001111100_0000100000000000"; -- 0.2831425666809082
	pesos_i(2106) := b"0000000000000000_0000000000000000_0001101101001011_1000101000000000"; -- 0.1066213846206665
	pesos_i(2107) := b"0000000000000000_0000000000000000_0010010110111100_1111101111000000"; -- 0.1474149078130722
	pesos_i(2108) := b"0000000000000000_0000000000000000_0001101110011100_0001101000000000"; -- 0.10785067081451416
	pesos_i(2109) := b"1111111111111111_1111111111111111_1100111001110011_1101010010000000"; -- -0.19354507327079773
	pesos_i(2110) := b"0000000000000000_0000000000000000_0010101001110110_0111111001000000"; -- 0.1658705621957779
	pesos_i(2111) := b"0000000000000000_0000000000000000_0000010001101101_0100100110011000"; -- 0.01729259453713894
	pesos_i(2112) := b"1111111111111111_1111111111111111_1111101111001001_0110001001110000"; -- -0.016458366066217422
	pesos_i(2113) := b"1111111111111111_1111111111111111_1110111110100111_1011001001000000"; -- -0.06384740769863129
	pesos_i(2114) := b"1111111111111111_1111111111111111_1100101000110101_0111001000000000"; -- -0.2101219892501831
	pesos_i(2115) := b"1111111111111111_1111111111111111_1110100000101011_0111011010000000"; -- -0.09308680891990662
	pesos_i(2116) := b"1111111111111111_1111111111111111_1111010011101110_0100101101010000"; -- -0.04323891922831535
	pesos_i(2117) := b"0000000000000000_0000000000000000_0011111111111100_0011000110000000"; -- 0.24994191527366638
	pesos_i(2118) := b"1111111111111111_1111111111111111_1110110110010100_0101100111100000"; -- -0.07195509225130081
	pesos_i(2119) := b"0000000000000000_0000000000000000_0010101101111001_1110010001000000"; -- 0.16982866823673248
	pesos_i(2120) := b"0000000000000000_0000000000000000_0100110101011101_1101111100000000"; -- 0.3022136092185974
	pesos_i(2121) := b"0000000000000000_0000000000000000_0000010000000010_0111001101100000"; -- 0.01566239446401596
	pesos_i(2122) := b"1111111111111111_1111111111111111_1101010100001110_1010011100000000"; -- -0.1677451729774475
	pesos_i(2123) := b"0000000000000000_0000000000000000_0010011111101110_1100001001000000"; -- 0.15598691999912262
	pesos_i(2124) := b"1111111111111111_1111111111111111_1110010001001100_0011011111000000"; -- -0.10821200907230377
	pesos_i(2125) := b"0000000000000000_0000000000000000_0110011100100100_0010101000000000"; -- 0.40289556980133057
	pesos_i(2126) := b"1111111111111111_1111111111111111_1001010101101101_0110001000000000"; -- -0.4162997007369995
	pesos_i(2127) := b"0000000000000000_0000000000000000_0000011010000011_1100001101111000"; -- 0.02544805221259594
	pesos_i(2128) := b"1111111111111111_1111111111111111_1101101000110110_0001101001000000"; -- -0.14761196076869965
	pesos_i(2129) := b"1111111111111111_1111111111111111_1110100000110100_1101001000000000"; -- -0.09294402599334717
	pesos_i(2130) := b"0000000000000000_0000000000000000_0001010101010101_0111110000000000"; -- 0.08333563804626465
	pesos_i(2131) := b"1111111111111111_1111111111111111_1110001110000101_0101011010100000"; -- -0.11124666780233383
	pesos_i(2132) := b"1111111111111111_1111111111111111_1111001010011000_1000111011110000"; -- -0.05235964432358742
	pesos_i(2133) := b"1111111111111111_1111111111111111_1110110110000011_1101010111100000"; -- -0.07220710068941116
	pesos_i(2134) := b"0000000000000000_0000000000000000_0000011010011011_0000110011010000"; -- 0.025803375989198685
	pesos_i(2135) := b"0000000000000000_0000000000000000_0010101010100100_0011000001000000"; -- 0.1665678173303604
	pesos_i(2136) := b"0000000000000000_0000000000000000_0010000101010100_1001101111000000"; -- 0.13019727170467377
	pesos_i(2137) := b"0000000000000000_0000000000000000_0010101101110010_1110100001000000"; -- 0.16972209513187408
	pesos_i(2138) := b"0000000000000000_0000000000000000_0001010110111000_0100000101000000"; -- 0.0848427563905716
	pesos_i(2139) := b"0000000000000000_0000000000000000_0001001100000010_1100001110100000"; -- 0.07426092773675919
	pesos_i(2140) := b"1111111111111111_1111111111111111_1010011001010000_0101100000000000"; -- -0.35033655166625977
	pesos_i(2141) := b"0000000000000000_0000000000000000_0001000000100011_1101111110100000"; -- 0.0630473867058754
	pesos_i(2142) := b"0000000000000000_0000000000000000_0010001110001101_0011010011000000"; -- 0.1388733834028244
	pesos_i(2143) := b"0000000000000000_0000000000000000_0100011000010000_0000011000000000"; -- 0.27368199825286865
	pesos_i(2144) := b"1111111111111111_1111111111111111_1101011001110101_1001011010000000"; -- -0.1622682511806488
	pesos_i(2145) := b"1111111111111111_1111111111111111_1111100010011111_0010011111000000"; -- -0.028821483254432678
	pesos_i(2146) := b"0000000000000000_0000000000000000_0011000101110000_1101010011000000"; -- 0.19312791526317596
	pesos_i(2147) := b"0000000000000000_0000000000000000_0000011110111111_0010101110111000"; -- 0.030260784551501274
	pesos_i(2148) := b"0000000000000000_0000000000000000_0010010111111000_0101110011000000"; -- 0.14832095801830292
	pesos_i(2149) := b"0000000000000000_0000000000000000_0001010101110111_0101001011100000"; -- 0.08385198563337326
	pesos_i(2150) := b"1111111111111111_1111111111111111_1110011010110101_0001110100100000"; -- -0.09879892319440842
	pesos_i(2151) := b"0000000000000000_0000000000000000_0000001101111011_0000000010011000"; -- 0.013595616444945335
	pesos_i(2152) := b"1111111111111111_1111111111111111_1100100010011110_0100000010000000"; -- -0.216335266828537
	pesos_i(2153) := b"0000000000000000_0000000000000000_0000010010010110_0000010101011000"; -- 0.01791413687169552
	pesos_i(2154) := b"1111111111111111_1111111111111111_1100110111010110_1111011011000000"; -- -0.19593866169452667
	pesos_i(2155) := b"0000000000000000_0000000000000000_0011100110111000_1000100010000000"; -- 0.22547200322151184
	pesos_i(2156) := b"0000000000000000_0000000000000000_0000110100100000_0010110000100000"; -- 0.051272161304950714
	pesos_i(2157) := b"1111111111111111_1111111111111111_1110000011110001_0011101110100000"; -- -0.12131907790899277
	pesos_i(2158) := b"1111111111111111_1111111111111111_1110100010010011_1111001000000000"; -- -0.09149253368377686
	pesos_i(2159) := b"1111111111111111_1111111111111111_1110110110011111_0001100111100000"; -- -0.07179106026887894
	pesos_i(2160) := b"1111111111111111_1111111111111111_1101100000010110_0001011010000000"; -- -0.15591296553611755
	pesos_i(2161) := b"1111111111111111_1111111111111111_1100000101001110_1000001110000000"; -- -0.24489572644233704
	pesos_i(2162) := b"0000000000000000_0000000000000000_0000010011010100_0001111111010000"; -- 0.018861759454011917
	pesos_i(2163) := b"0000000000000000_0000000000000000_0000111011001001_1001010000000000"; -- 0.05776333808898926
	pesos_i(2164) := b"1111111111111111_1111111111111111_1111010000101101_1011000110110000"; -- -0.04617776349186897
	pesos_i(2165) := b"1111111111111111_1111111111111111_1100110100010001_1001100101000000"; -- -0.19895021617412567
	pesos_i(2166) := b"0000000000000000_0000000000000000_0100010010010000_0111010110000000"; -- 0.2678292691707611
	pesos_i(2167) := b"0000000000000000_0000000000000000_0001010011001000_0111001100000000"; -- 0.08118361234664917
	pesos_i(2168) := b"0000000000000000_0000000000000000_0011110011001010_1100011011000000"; -- 0.2374691218137741
	pesos_i(2169) := b"0000000000000000_0000000000000000_0100111011110011_1011000000000000"; -- 0.30840587615966797
	pesos_i(2170) := b"1111111111111111_1111111111111111_1100001000101101_0001011010000000"; -- -0.24149951338768005
	pesos_i(2171) := b"1111111111111111_1111111111111111_1100111110001101_0111100000000000"; -- -0.18924760818481445
	pesos_i(2172) := b"1111111111111111_1111111111111111_1110111000000001_0101100111100000"; -- -0.07029188424348831
	pesos_i(2173) := b"0000000000000000_0000000000000000_0010110110101000_1110111101000000"; -- 0.1783589869737625
	pesos_i(2174) := b"1111111111111111_1111111111111111_1110101111001110_0010111011100000"; -- -0.07888514548540115
	pesos_i(2175) := b"1111111111111111_1111111111111111_1110100100011010_0010110000000000"; -- -0.08944439888000488
	pesos_i(2176) := b"1111111111111111_1111111111111111_1111110101011000_1110001011110000"; -- -0.010362450033426285
	pesos_i(2177) := b"1111111111111111_1111111111111111_1111111111000000_0101110101111111"; -- -0.0009709896985441446
	pesos_i(2178) := b"0000000000000000_0000000000000000_0001111111001011_0111101101000000"; -- 0.12419863045215607
	pesos_i(2179) := b"0000000000000000_0000000000000000_0000011101101011_0000101101111000"; -- 0.028977124020457268
	pesos_i(2180) := b"0000000000000000_0000000000000000_0001000001100011_1001011111000000"; -- 0.06401966512203217
	pesos_i(2181) := b"1111111111111111_1111111111111111_1011001010001010_1101100010000000"; -- -0.30256888270378113
	pesos_i(2182) := b"1111111111111111_1111111111111111_1111100111101001_0010011000000000"; -- -0.023786187171936035
	pesos_i(2183) := b"0000000000000000_0000000000000000_0000101101111011_0001110000000000"; -- 0.04484724998474121
	pesos_i(2184) := b"0000000000000000_0000000000000000_0011100001101110_0010000110000000"; -- 0.22043046355247498
	pesos_i(2185) := b"1111111111111111_1111111111111111_1100110101001100_0100011110000000"; -- -0.19805482029914856
	pesos_i(2186) := b"0000000000000000_0000000000000000_0000000001011000_1001000111101100"; -- 0.0013514709426090121
	pesos_i(2187) := b"0000000000000000_0000000000000000_0101001001101011_0000100010000000"; -- 0.3219456970691681
	pesos_i(2188) := b"0000000000000000_0000000000000000_0001010100010001_0101101111100000"; -- 0.08229612559080124
	pesos_i(2189) := b"1111111111111111_1111111111111111_1110101111101010_1011010001100000"; -- -0.07844994217157364
	pesos_i(2190) := b"1111111111111111_1111111111111111_1111101010011001_1000111000001000"; -- -0.021094439551234245
	pesos_i(2191) := b"0000000000000000_0000000000000000_0000101111000000_1001101100110000"; -- 0.04590768739581108
	pesos_i(2192) := b"1111111111111111_1111111111111111_1000110011100101_1000011000000000"; -- -0.4496227502822876
	pesos_i(2193) := b"1111111111111111_1111111111111111_1111110100111110_1010110111011000"; -- -0.010762343183159828
	pesos_i(2194) := b"1111111111111111_1111111111111111_1100110101110010_1100111001000000"; -- -0.19746695458889008
	pesos_i(2195) := b"1111111111111111_1111111111111111_1110001101100000_1011110101000000"; -- -0.11180512607097626
	pesos_i(2196) := b"0000000000000000_0000000000000000_0001110011011011_0011001110100000"; -- 0.11271975189447403
	pesos_i(2197) := b"0000000000000000_0000000000000000_0000011010000101_1110101111000000"; -- 0.0254809707403183
	pesos_i(2198) := b"0000000000000000_0000000000000000_0001100100110101_1100000000000000"; -- 0.09847640991210938
	pesos_i(2199) := b"0000000000000000_0000000000000000_0010000001111110_0011010010000000"; -- 0.1269257366657257
	pesos_i(2200) := b"1111111111111111_1111111111111111_1100111001001010_0000110010000000"; -- -0.1941826045513153
	pesos_i(2201) := b"1111111111111111_1111111111111111_1111111101011000_0011100100001100"; -- -0.002560076303780079
	pesos_i(2202) := b"0000000000000000_0000000000000000_0000110010011000_1111111001100000"; -- 0.04920949786901474
	pesos_i(2203) := b"1111111111111111_1111111111111111_1110110111001000_1110111010100000"; -- -0.07115276902914047
	pesos_i(2204) := b"0000000000000000_0000000000000000_0010100101001101_1011010001000000"; -- 0.16134192049503326
	pesos_i(2205) := b"0000000000000000_0000000000000000_0001101011001110_1101100100000000"; -- 0.10471874475479126
	pesos_i(2206) := b"0000000000000000_0000000000000000_0001011001001001_0000000001100000"; -- 0.08705141395330429
	pesos_i(2207) := b"0000000000000000_0000000000000000_0010101100001111_1000011111000000"; -- 0.16820572316646576
	pesos_i(2208) := b"1111111111111111_1111111111111111_1011110100010110_1110000100000000"; -- -0.26136964559555054
	pesos_i(2209) := b"1111111111111111_1111111111111111_1111110101110100_1101010000000000"; -- -0.009936094284057617
	pesos_i(2210) := b"0000000000000000_0000000000000000_0001111111111011_1101011010100000"; -- 0.12493649870157242
	pesos_i(2211) := b"1111111111111111_1111111111111111_1100111000001111_0011111110000000"; -- -0.19507983326911926
	pesos_i(2212) := b"1111111111111111_1111111111111111_1101010111100010_0011010011000000"; -- -0.1645171195268631
	pesos_i(2213) := b"0000000000000000_0000000000000000_0000110110010011_1010101100010000"; -- 0.05303448811173439
	pesos_i(2214) := b"1111111111111111_1111111111111111_1101000000101101_1110010000000000"; -- -0.1867997646331787
	pesos_i(2215) := b"1111111111111111_1111111111111111_1110111110111000_0101001000000000"; -- -0.06359374523162842
	pesos_i(2216) := b"1111111111111111_1111111111111111_1111000001011101_0111000101010000"; -- -0.06107417866587639
	pesos_i(2217) := b"0000000000000000_0000000000000000_0001000110111101_0001001000100000"; -- 0.06929124146699905
	pesos_i(2218) := b"0000000000000000_0000000000000000_0001000000101001_1001001111000000"; -- 0.06313441693782806
	pesos_i(2219) := b"1111111111111111_1111111111111111_1100010011101110_1100011100000000"; -- -0.2307315468788147
	pesos_i(2220) := b"0000000000000000_0000000000000000_0001011010100000_0101010111000000"; -- 0.08838401734828949
	pesos_i(2221) := b"0000000000000000_0000000000000000_0000101110001110_0010011011000000"; -- 0.045137807726860046
	pesos_i(2222) := b"0000000000000000_0000000000000000_0100001001110011_1100001000000000"; -- 0.2595788240432739
	pesos_i(2223) := b"0000000000000000_0000000000000000_0011000010000001_1001000110000000"; -- 0.18947705626487732
	pesos_i(2224) := b"0000000000000000_0000000000000000_0001101001011110_0010010001000000"; -- 0.10299898684024811
	pesos_i(2225) := b"1111111111111111_1111111111111111_1111001000011001_1011110100100000"; -- -0.054294757544994354
	pesos_i(2226) := b"1111111111111111_1111111111111111_1110111001010001_0001010111000000"; -- -0.06907524168491364
	pesos_i(2227) := b"0000000000000000_0000000000000000_0000000001001100_1001101000001100"; -- 0.001168849878013134
	pesos_i(2228) := b"0000000000000000_0000000000000000_0000011110010010_1101111011001000"; -- 0.029584812000393867
	pesos_i(2229) := b"0000000000000000_0000000000000000_0000000011111111_0011111011101110"; -- 0.003894742112606764
	pesos_i(2230) := b"0000000000000000_0000000000000000_0010010000001010_0000010111000000"; -- 0.14077793061733246
	pesos_i(2231) := b"0000000000000000_0000000000000000_0011001111000111_0101100101000000"; -- 0.2022605687379837
	pesos_i(2232) := b"1111111111111111_1111111111111111_1101000110001111_0100010101000000"; -- -0.1814076155424118
	pesos_i(2233) := b"0000000000000000_0000000000000000_0100101101011010_1101000110000000"; -- 0.29435452818870544
	pesos_i(2234) := b"1111111111111111_1111111111111111_1110111101100100_1000100000100000"; -- -0.06487225741147995
	pesos_i(2235) := b"0000000000000000_0000000000000000_0000111001001101_0101111101010000"; -- 0.055868107825517654
	pesos_i(2236) := b"0000000000000000_0000000000000000_0100111011111101_1101101110000000"; -- 0.3085610568523407
	pesos_i(2237) := b"1111111111111111_1111111111111111_1000111000101110_0111001010000000"; -- -0.4446037709712982
	pesos_i(2238) := b"0000000000000000_0000000000000000_0001100111101110_0100010011000000"; -- 0.10129193961620331
	pesos_i(2239) := b"1111111111111111_1111111111111111_1111000011001011_1010011110000000"; -- -0.05939248204231262
	pesos_i(2240) := b"1111111111111111_1111111111111111_1101011101010011_0000010000000000"; -- -0.1588895320892334
	pesos_i(2241) := b"1111111111111111_1111111111111111_1101110010100001_0010111111000000"; -- -0.13816548883914948
	pesos_i(2242) := b"0000000000000000_0000000000000000_0000001100110101_1010111110100000"; -- 0.012537933886051178
	pesos_i(2243) := b"0000000000000000_0000000000000000_0001100001100000_1100110101000000"; -- 0.09522707760334015
	pesos_i(2244) := b"0000000000000000_0000000000000000_0010101001110110_1111100100000000"; -- 0.16587787866592407
	pesos_i(2245) := b"0000000000000000_0000000000000000_0100001110000111_0110011000000000"; -- 0.2637847661972046
	pesos_i(2246) := b"1111111111111111_1111111111111111_1110010001011001_0000010111000000"; -- -0.10801662504673004
	pesos_i(2247) := b"0000000000000000_0000000000000000_0001111011010000_1000110011000000"; -- 0.12036971747875214
	pesos_i(2248) := b"1111111111111111_1111111111111111_1011110011000101_1001100110000000"; -- -0.2626098692417145
	pesos_i(2249) := b"1111111111111111_1111111111111111_1110001010011001_0010011101100000"; -- -0.11485055834054947
	pesos_i(2250) := b"0000000000000000_0000000000000000_0000100001010111_0100000010010000"; -- 0.03258136287331581
	pesos_i(2251) := b"1111111111111111_1111111111111111_1111100100011110_1100111100111000"; -- -0.02687363512814045
	pesos_i(2252) := b"1111111111111111_1111111111111111_1100110001010110_1001011000000000"; -- -0.2018038034439087
	pesos_i(2253) := b"0000000000000000_0000000000000000_0110010101000011_0000001110000000"; -- 0.3955537974834442
	pesos_i(2254) := b"1111111111111111_1111111111111111_1100110010111100_1010011001000000"; -- -0.2002464383840561
	pesos_i(2255) := b"1111111111111111_1111111111111111_1110010101100000_1111100100000000"; -- -0.10398906469345093
	pesos_i(2256) := b"0000000000000000_0000000000000000_0000010111001101_0101110101000000"; -- 0.022664859890937805
	pesos_i(2257) := b"1111111111111111_1111111111111111_1110110111001101_1101111010000000"; -- -0.07107743620872498
	pesos_i(2258) := b"1111111111111111_1111111111111111_1110011000110000_1010010111100000"; -- -0.10082019120454788
	pesos_i(2259) := b"0000000000000000_0000000000000000_0000111000101011_1010111100110000"; -- 0.05535406991839409
	pesos_i(2260) := b"0000000000000000_0000000000000000_0010100101001010_1000001100000000"; -- 0.16129320859909058
	pesos_i(2261) := b"0000000000000000_0000000000000000_0011010010010111_1011001000000000"; -- 0.20543968677520752
	pesos_i(2262) := b"1111111111111111_1111111111111111_1110000000100101_0110010011100000"; -- -0.12442941218614578
	pesos_i(2263) := b"0000000000000000_0000000000000000_0100001111101111_1010111000000000"; -- 0.2653759717941284
	pesos_i(2264) := b"0000000000000000_0000000000000000_0001011010000110_1000010110000000"; -- 0.08799013495445251
	pesos_i(2265) := b"1111111111111111_1111111111111111_1011111111111110_0010000000000000"; -- -0.2500286102294922
	pesos_i(2266) := b"0000000000000000_0000000000000000_0011011101110011_1111110011000000"; -- 0.21661357581615448
	pesos_i(2267) := b"1111111111111111_1111111111111111_1111101001110100_1111101111000000"; -- -0.021652474999427795
	pesos_i(2268) := b"0000000000000000_0000000000000000_0001011100110010_1110011001000000"; -- 0.09062041342258453
	pesos_i(2269) := b"0000000000000000_0000000000000000_0000101001011011_0101100111110000"; -- 0.04045641049742699
	pesos_i(2270) := b"0000000000000000_0000000000000000_0001101000010011_1111001111100000"; -- 0.1018669530749321
	pesos_i(2271) := b"0000000000000000_0000000000000000_0000010010010000_0001011111011000"; -- 0.017823686823248863
	pesos_i(2272) := b"1111111111111111_1111111111111111_1101011000100000_0011111111000000"; -- -0.16357041895389557
	pesos_i(2273) := b"1111111111111111_1111111111111111_1111100000110011_1001011110001000"; -- -0.03046276979148388
	pesos_i(2274) := b"1111111111111111_1111111111111111_1111000000011110_0001001000010000"; -- -0.062041159719228745
	pesos_i(2275) := b"1111111111111111_1111111111111111_1111101101001011_0111001100001000"; -- -0.01837998442351818
	pesos_i(2276) := b"0000000000000000_0000000000000000_0001000000100011_1110010101000000"; -- 0.06304772198200226
	pesos_i(2277) := b"0000000000000000_0000000000000000_0001101100001001_0101011100000000"; -- 0.10561126470565796
	pesos_i(2278) := b"1111111111111111_1111111111111111_1010010011101000_1011000000000000"; -- -0.35582447052001953
	pesos_i(2279) := b"1111111111111111_1111111111111111_1110010001010101_1111110111100000"; -- -0.10806287080049515
	pesos_i(2280) := b"1111111111111111_1111111111111111_1111100111110011_1110001011110000"; -- -0.023622337728738785
	pesos_i(2281) := b"0000000000000000_0000000000000000_0001010011110011_0110011011100000"; -- 0.08183901757001877
	pesos_i(2282) := b"1111111111111111_1111111111111111_1111100011010101_1101110000111000"; -- -0.02798675186932087
	pesos_i(2283) := b"0000000000000000_0000000000000000_0000101010010010_1111000110010000"; -- 0.041304681450128555
	pesos_i(2284) := b"1111111111111111_1111111111111111_1110011000101011_1000110100100000"; -- -0.10089796036481857
	pesos_i(2285) := b"1111111111111111_1111111111111111_1100110111101100_1111011010000000"; -- -0.19560298323631287
	pesos_i(2286) := b"1111111111111111_1111111111111111_1110010101011111_1000011111000000"; -- -0.10401107370853424
	pesos_i(2287) := b"0000000000000000_0000000000000000_0000000101000100_1010110101011000"; -- 0.004954179748892784
	pesos_i(2288) := b"0000000000000000_0000000000000000_0010000101010100_1101101011000000"; -- 0.13020102679729462
	pesos_i(2289) := b"1111111111111111_1111111111111111_1111100111101001_0110110000100000"; -- -0.02378200739622116
	pesos_i(2290) := b"1111111111111111_1111111111111111_1111110010101111_1000001101111100"; -- -0.01294687483459711
	pesos_i(2291) := b"0000000000000000_0000000000000000_0100011111010001_0010101110000000"; -- 0.28053542971611023
	pesos_i(2292) := b"1111111111111111_1111111111111111_1111110110000110_0010000001110100"; -- -0.009672137908637524
	pesos_i(2293) := b"1111111111111111_1111111111111111_1011111100101110_1110100110000000"; -- -0.25319042801856995
	pesos_i(2294) := b"0000000000000000_0000000000000000_0000110001110100_1100011111100000"; -- 0.04865693300962448
	pesos_i(2295) := b"0000000000000000_0000000000000000_0011110000001110_1111001001000000"; -- 0.23460306227207184
	pesos_i(2296) := b"1111111111111111_1111111111111111_1100011010001001_0001100000000000"; -- -0.2244706153869629
	pesos_i(2297) := b"0000000000000000_0000000000000000_0100001111101110_0000100100000000"; -- 0.265350878238678
	pesos_i(2298) := b"1111111111111111_1111111111111111_1101001001111011_0011110100000000"; -- -0.1778070330619812
	pesos_i(2299) := b"0000000000000000_0000000000000000_0000101001111000_0101100100110000"; -- 0.040898870676755905
	pesos_i(2300) := b"1111111111111111_1111111111111111_1011001010110001_0101000100000000"; -- -0.3019818663597107
	pesos_i(2301) := b"1111111111111111_1111111111111111_1111000100110010_1010111011000000"; -- -0.0578203946352005
	pesos_i(2302) := b"1111111111111111_1111111111111111_1101000101101101_1101000011000000"; -- -0.18191809952259064
	pesos_i(2303) := b"1111111111111111_1111111111111111_1101000000111100_1000111000000000"; -- -0.1865760087966919
	pesos_i(2304) := b"0000000000000000_0000000000000000_0001110010110010_0101011110100000"; -- 0.11209628731012344
	pesos_i(2305) := b"0000000000000000_0000000000000000_0010101000111101_0001000011000000"; -- 0.1649942845106125
	pesos_i(2306) := b"0000000000000000_0000000000000000_0011101000110110_1011111011000000"; -- 0.2273978441953659
	pesos_i(2307) := b"0000000000000000_0000000000000000_0011111111101100_0000110001000000"; -- 0.2496955543756485
	pesos_i(2308) := b"0000000000000000_0000000000000000_0011001110000001_0000001110000000"; -- 0.2011873424053192
	pesos_i(2309) := b"1111111111111111_1111111111111111_0100111101000101_0111111100000000"; -- -0.690345823764801
	pesos_i(2310) := b"0000000000000000_0000000000000000_0010010011101100_1111110100000000"; -- 0.14424115419387817
	pesos_i(2311) := b"0000000000000000_0000000000000000_0000101011000010_1001010000110000"; -- 0.04203153774142265
	pesos_i(2312) := b"0000000000000000_0000000000000000_0011111000101010_0001111111000000"; -- 0.24283026158809662
	pesos_i(2313) := b"0000000000000000_0000000000000000_0011000000100101_1111101001000000"; -- 0.18807949125766754
	pesos_i(2314) := b"0000000000000000_0000000000000000_0010010010110010_0000111011000000"; -- 0.14334194362163544
	pesos_i(2315) := b"0000000000000000_0000000000000000_0011000101001101_1001011011000000"; -- 0.1925901621580124
	pesos_i(2316) := b"0000000000000000_0000000000000000_0011001011100001_1011010000000000"; -- 0.19875645637512207
	pesos_i(2317) := b"1111111111111111_1111111111111111_1100100111000001_1111001001000000"; -- -0.21188436448574066
	pesos_i(2318) := b"1111111111111111_1111111111111111_0101111111010100_0101111000000000"; -- -0.6256657838821411
	pesos_i(2319) := b"1111111111111111_1111111111111111_1110100011100110_1111111000100000"; -- -0.09022533148527145
	pesos_i(2320) := b"1111111111111111_1111111111111111_1110001001101000_1011100111000000"; -- -0.11558951437473297
	pesos_i(2321) := b"0000000000000000_0000000000000000_0010010001111010_0001100000000000"; -- 0.1424880027770996
	pesos_i(2322) := b"1111111111111111_1111111111111111_1110100110000111_0111010111000000"; -- -0.0877767950296402
	pesos_i(2323) := b"1111111111111111_1111111111111111_1101101010100011_0011011111000000"; -- -0.14594699442386627
	pesos_i(2324) := b"0000000000000000_0000000000000000_0101001001000110_1100010100000000"; -- 0.32139235734939575
	pesos_i(2325) := b"1111111111111111_1111111111111111_1110111001001110_1110010000100000"; -- -0.06910871714353561
	pesos_i(2326) := b"0000000000000000_0000000000000000_0011000010101111_0010000001000000"; -- 0.1901722103357315
	pesos_i(2327) := b"0000000000000000_0000000000000000_0001101101000011_0110000000100000"; -- 0.10649681836366653
	pesos_i(2328) := b"1111111111111111_1111111111111111_1110011101000101_0100111000100000"; -- -0.09659873694181442
	pesos_i(2329) := b"0000000000000000_0000000000000000_0101100001010111_0100000000000000"; -- 0.3450813293457031
	pesos_i(2330) := b"0000000000000000_0000000000000000_0000100111101000_0011001000110000"; -- 0.038699280470609665
	pesos_i(2331) := b"0000000000000000_0000000000000000_0000110110100000_1110001101100000"; -- 0.053236208856105804
	pesos_i(2332) := b"1111111111111111_1111111111111111_1011100110111100_1101110010000000"; -- -0.274461954832077
	pesos_i(2333) := b"0000000000000000_0000000000000000_0101010001000000_1010001000000000"; -- 0.3291112184524536
	pesos_i(2334) := b"0000000000000000_0000000000000000_0011010000000000_0100000000000000"; -- 0.20312881469726562
	pesos_i(2335) := b"0000000000000000_0000000000000000_0011100000011110_0010100011000000"; -- 0.2192101925611496
	pesos_i(2336) := b"1111111111111111_1111111111111111_1100110011110000_0001101001000000"; -- -0.19946132600307465
	pesos_i(2337) := b"1111111111111111_1111111111111111_1111100000100111_0111010011010000"; -- -0.030647944658994675
	pesos_i(2338) := b"0000000000000000_0000000000000000_0100111000110110_1110000110000000"; -- 0.30552491545677185
	pesos_i(2339) := b"0000000000000000_0000000000000000_0011011011001001_0000001000000000"; -- 0.21400463581085205
	pesos_i(2340) := b"1111111111111111_1111111111111111_1001000110100110_1111001110000000"; -- -0.4310462772846222
	pesos_i(2341) := b"0000000000000000_0000000000000000_0000011110000001_0101110010110000"; -- 0.02931765839457512
	pesos_i(2342) := b"0000000000000000_0000000000000000_0010110111101111_0001011011000000"; -- 0.17942945659160614
	pesos_i(2343) := b"0000000000000000_0000000000000000_0001111111101001_1100111000000000"; -- 0.12466132640838623
	pesos_i(2344) := b"0000000000000000_0000000000000000_0001101000110001_1011101100100000"; -- 0.1023213341832161
	pesos_i(2345) := b"1111111111111111_1111111111111111_1101101001100011_1110001011000000"; -- -0.14691336452960968
	pesos_i(2346) := b"1111111111111111_1111111111111111_1110011001100100_1010111001100000"; -- -0.10002622753381729
	pesos_i(2347) := b"1111111111111111_1111111111111111_1011101101011000_0001000110000000"; -- -0.26818743348121643
	pesos_i(2348) := b"1111111111111111_1111111111111111_1101001000101010_0100101011000000"; -- -0.17904217541217804
	pesos_i(2349) := b"0000000000000000_0000000000000000_0001011111101100_0100101100000000"; -- 0.09344929456710815
	pesos_i(2350) := b"0000000000000000_0000000000000000_0011101000010010_1110001011000000"; -- 0.22685067355632782
	pesos_i(2351) := b"0000000000000000_0000000000000000_0101001110011010_0011111110000000"; -- 0.32657238841056824
	pesos_i(2352) := b"0000000000000000_0000000000000000_0000000100101001_0011100000001100"; -- 0.004535201005637646
	pesos_i(2353) := b"0000000000000000_0000000000000000_0000100011000000_0001110101110000"; -- 0.034181442111730576
	pesos_i(2354) := b"1111111111111111_1111111111111111_1110110111001001_1010101100000000"; -- -0.07114154100418091
	pesos_i(2355) := b"0000000000000000_0000000000000000_0010000100110010_0000010100000000"; -- 0.12966948747634888
	pesos_i(2356) := b"0000000000000000_0000000000000000_0101101011100100_0011101100000000"; -- 0.35504502058029175
	pesos_i(2357) := b"0000000000000000_0000000000000000_0001111111100101_0010010111100000"; -- 0.12459027022123337
	pesos_i(2358) := b"0000000000000000_0000000000000000_0011011010111001_0111011101000000"; -- 0.21376748383045197
	pesos_i(2359) := b"0000000000000000_0000000000000000_0101100111000101_1101100100000000"; -- 0.35067516565322876
	pesos_i(2360) := b"1111111111111111_1111111111111111_1111100011001100_1100000001100000"; -- -0.028125740587711334
	pesos_i(2361) := b"0000000000000000_0000000000000000_0010111010111100_0111111001000000"; -- 0.1825636774301529
	pesos_i(2362) := b"0000000000000000_0000000000000000_0001110101011001_0010100010100000"; -- 0.1146417036652565
	pesos_i(2363) := b"1111111111111111_1111111111111111_1101000011001110_1100001100000000"; -- -0.1843450665473938
	pesos_i(2364) := b"1111111111111111_1111111111111111_1111110111101111_0001001111001000"; -- -0.008070720359683037
	pesos_i(2365) := b"1111111111111111_1111111111111111_1101010000111111_1111011110000000"; -- -0.1708989441394806
	pesos_i(2366) := b"0000000000000000_0000000000000000_0100110101101100_1101111100000000"; -- 0.3024424910545349
	pesos_i(2367) := b"0000000000000000_0000000000000000_0011101011111111_0110111011000000"; -- 0.23046009242534637
	pesos_i(2368) := b"1111111111111111_1111111111111111_1110111000001000_1110111010100000"; -- -0.07017620652914047
	pesos_i(2369) := b"1111111111111111_1111111111111111_1011100001001110_0111010010000000"; -- -0.28005287051200867
	pesos_i(2370) := b"1111111111111111_1111111111111111_1100010010000000_0001010111000000"; -- -0.23242057859897614
	pesos_i(2371) := b"0000000000000000_0000000000000000_0010000101111110_1001010100000000"; -- 0.13083773851394653
	pesos_i(2372) := b"0000000000000000_0000000000000000_0001000011111111_0111010110000000"; -- 0.06639799475669861
	pesos_i(2373) := b"0000000000000000_0000000000000000_0010111010011110_0111011010000000"; -- 0.18210545182228088
	pesos_i(2374) := b"1111111111111111_1111111111111111_0011111111110001_0111110000000000"; -- -0.7502214908599854
	pesos_i(2375) := b"0000000000000000_0000000000000000_0100010010101010_0101110010000000"; -- 0.2682245075702667
	pesos_i(2376) := b"1111111111111111_1111111111111111_0110010010010111_0101000000000000"; -- -0.6070661544799805
	pesos_i(2377) := b"0000000000000000_0000000000000000_0010000110010000_0101100011000000"; -- 0.13110880553722382
	pesos_i(2378) := b"1111111111111111_1111111111111111_1110101001011010_1111010100000000"; -- -0.08454960584640503
	pesos_i(2379) := b"1111111111111111_1111111111111111_1100011011111010_1010010100000000"; -- -0.22273796796798706
	pesos_i(2380) := b"0000000000000000_0000000000000000_0010001111001010_1010101001000000"; -- 0.139811173081398
	pesos_i(2381) := b"0000000000000000_0000000000000000_0001111000011011_1100011100100000"; -- 0.1176113560795784
	pesos_i(2382) := b"1111111111111111_1111111111111111_1100011110001011_1011111011000000"; -- -0.2205239087343216
	pesos_i(2383) := b"1111111111111111_1111111111111111_1011000001011001_0111011000000000"; -- -0.311134934425354
	pesos_i(2384) := b"1111111111111111_1111111111111111_1100111001010101_1100000000000000"; -- -0.19400405883789062
	pesos_i(2385) := b"0000000000000000_0000000000000000_0011011010011100_0000011011000000"; -- 0.21331827342510223
	pesos_i(2386) := b"1111111111111111_1111111111111111_1111000110101011_1110011111110000"; -- -0.05597067251801491
	pesos_i(2387) := b"1111111111111111_1111111111111111_1111010111000001_1110001001010000"; -- -0.04001031443476677
	pesos_i(2388) := b"0000000000000000_0000000000000000_0110000000001001_0001111100000000"; -- 0.37513917684555054
	pesos_i(2389) := b"0000000000000000_0000000000000000_0011001001011111_0101101110000000"; -- 0.19676753878593445
	pesos_i(2390) := b"1111111111111111_1111111111111111_1111110001001011_0110000101001100"; -- -0.01447479147464037
	pesos_i(2391) := b"0000000000000000_0000000000000000_0111000010101011_1010110000000000"; -- 0.44011950492858887
	pesos_i(2392) := b"0000000000000000_0000000000000000_0011111101010101_1001111100000000"; -- 0.2474002242088318
	pesos_i(2393) := b"0000000000000000_0000000000000000_0001000011110000_1000100011000000"; -- 0.06617026031017303
	pesos_i(2394) := b"1111111111111111_1111111111111111_1111000110111000_1110000110010000"; -- -0.05577268823981285
	pesos_i(2395) := b"1111111111111111_1111111111111111_1110100110010001_1100000110100000"; -- -0.08761968463659286
	pesos_i(2396) := b"0000000000000000_0000000000000000_0011000110011001_0101001010000000"; -- 0.19374576210975647
	pesos_i(2397) := b"0000000000000000_0000000000000000_0011101000011001_1100000000000000"; -- 0.22695541381835938
	pesos_i(2398) := b"1111111111111111_1111111111111111_1111111101010111_1000001000111001"; -- -0.002570973476395011
	pesos_i(2399) := b"1111111111111111_1111111111111111_1010010100010011_1011100000000000"; -- -0.35516786575317383
	pesos_i(2400) := b"1111111111111111_1111111111111111_1010100100001001_1011100000000000"; -- -0.33969545364379883
	pesos_i(2401) := b"1111111111111111_1111111111111111_1111111000111010_0001010110110000"; -- -0.006926197558641434
	pesos_i(2402) := b"0000000000000000_0000000000000000_0000111100100101_1001000001000000"; -- 0.05916692316532135
	pesos_i(2403) := b"0000000000000000_0000000000000000_0001001001100000_1010010001000000"; -- 0.07178713381290436
	pesos_i(2404) := b"1111111111111111_1111111111111111_1110100010010001_1101111011000000"; -- -0.09152419865131378
	pesos_i(2405) := b"0000000000000000_0000000000000000_0100100101001001_0000001100000000"; -- 0.2862703204154968
	pesos_i(2406) := b"1111111111111111_1111111111111111_1110111010110111_1000010100000000"; -- -0.06751221418380737
	pesos_i(2407) := b"0000000000000000_0000000000000000_0000100001110011_0111000001010000"; -- 0.033011455088853836
	pesos_i(2408) := b"0000000000000000_0000000000000000_0100100011110001_0010010000000000"; -- 0.2849295139312744
	pesos_i(2409) := b"1111111111111111_1111111111111111_1101101110001010_1100100111000000"; -- -0.14241351187229156
	pesos_i(2410) := b"0000000000000000_0000000000000000_0011001100000011_0100011001000000"; -- 0.19926871359348297
	pesos_i(2411) := b"1111111111111111_1111111111111111_1110111100101011_0000101011000000"; -- -0.06574948132038116
	pesos_i(2412) := b"1111111111111111_1111111111111111_1000101000110110_1001010110000000"; -- -0.4601046144962311
	pesos_i(2413) := b"1111111111111111_1111111111111111_1101010000000010_1010110001000000"; -- -0.17183421552181244
	pesos_i(2414) := b"0000000000000000_0000000000000000_0011100001001011_0010101000000000"; -- 0.21989691257476807
	pesos_i(2415) := b"0000000000000000_0000000000000000_0100000101001111_0011010010000000"; -- 0.2551148235797882
	pesos_i(2416) := b"1111111111111111_1111111111111111_1111100001110001_0100100011000000"; -- -0.02952142059803009
	pesos_i(2417) := b"0000000000000000_0000000000000000_0001111011010101_1100000011100000"; -- 0.12044911831617355
	pesos_i(2418) := b"0000000000000000_0000000000000000_0011110101001111_1101011000000000"; -- 0.23949944972991943
	pesos_i(2419) := b"0000000000000000_0000000000000000_0100001010010010_1010111100000000"; -- 0.2600507140159607
	pesos_i(2420) := b"0000000000000000_0000000000000000_0000111000010001_0010011000000000"; -- 0.054949164390563965
	pesos_i(2421) := b"1111111111111111_1111111111111111_1101000111000101_0110000000000000"; -- -0.18058204650878906
	pesos_i(2422) := b"1111111111111111_1111111111111111_1101100110010010_0101111111000000"; -- -0.15011025965213776
	pesos_i(2423) := b"1111111111111111_1111111111111111_1011110010101111_0100110100000000"; -- -0.2629501223564148
	pesos_i(2424) := b"1111111111111111_1111111111111111_1011001101101000_0110101000000000"; -- -0.2991880178451538
	pesos_i(2425) := b"0000000000000000_0000000000000000_0010101100000011_0110110010000000"; -- 0.16802099347114563
	pesos_i(2426) := b"1111111111111111_1111111111111111_1111011110011111_0100100001100000"; -- -0.03272578865289688
	pesos_i(2427) := b"0000000000000000_0000000000000000_0010100011111111_0101100000000000"; -- 0.16014623641967773
	pesos_i(2428) := b"0000000000000000_0000000000000000_0000011110101000_0110011111111000"; -- 0.02991342358291149
	pesos_i(2429) := b"1111111111111111_1111111111111111_1101010111001010_0000101011000000"; -- -0.16488583385944366
	pesos_i(2430) := b"0000000000000000_0000000000000000_0000010111001011_0010001000100000"; -- 0.02263081818819046
	pesos_i(2431) := b"1111111111111111_1111111111111111_1110100000111101_0010010010000000"; -- -0.0928170382976532
	pesos_i(2432) := b"1111111111111111_1111111111111111_1101101010000001_1000111000000000"; -- -0.1464606523513794
	pesos_i(2433) := b"0000000000000000_0000000000000000_1010010011000111_0101101000000000"; -- 0.6436668634414673
	pesos_i(2434) := b"0000000000000000_0000000000000000_0001100110000101_0101100101100000"; -- 0.0996909961104393
	pesos_i(2435) := b"0000000000000000_0000000000000000_0010000001111110_0010001110000000"; -- 0.12692472338676453
	pesos_i(2436) := b"1111111111111111_1111111111111111_1110011111001100_1100110110100000"; -- -0.09453120082616806
	pesos_i(2437) := b"1111111111111111_1111111111111111_1010011101011001_0011111100000000"; -- -0.34629446268081665
	pesos_i(2438) := b"1111111111111111_1111111111111111_1101010110000111_1010010100000000"; -- -0.16589897871017456
	pesos_i(2439) := b"1111111111111111_1111111111111111_1110011010001101_1010110101000000"; -- -0.09940068423748016
	pesos_i(2440) := b"0000000000000000_0000000000000000_0000111001000001_1001100110010000"; -- 0.05568847432732582
	pesos_i(2441) := b"0000000000000000_0000000000000000_0110100111110011_1001111100000000"; -- 0.4138736128807068
	pesos_i(2442) := b"1111111111111111_1111111111111111_1101101111000101_1101100000000000"; -- -0.14151239395141602
	pesos_i(2443) := b"0000000000000000_0000000000000000_0011100101101010_0000010100000000"; -- 0.22427397966384888
	pesos_i(2444) := b"0000000000000000_0000000000000000_0011011000001100_1010000010000000"; -- 0.21113017201423645
	pesos_i(2445) := b"1111111111111111_1111111111111111_1001100100101001_0110001010000000"; -- -0.4017122685909271
	pesos_i(2446) := b"1111111111111111_1111111111111111_1001111001110110_1001100100000000"; -- -0.38100284337997437
	pesos_i(2447) := b"1111111111111111_1111111111111111_1101110010110100_0000001000000000"; -- -0.13787829875946045
	pesos_i(2448) := b"0000000000000000_0000000000000000_0000101101111010_1100111100000000"; -- 0.044842660427093506
	pesos_i(2449) := b"1111111111111111_1111111111111111_1111011010111100_0000001101010000"; -- -0.03619365021586418
	pesos_i(2450) := b"0000000000000000_0000000000000000_0010000100100111_1101101001000000"; -- 0.12951435148715973
	pesos_i(2451) := b"1111111111111111_1111111111111111_1110110001011101_1110000000000000"; -- -0.07669258117675781
	pesos_i(2452) := b"1111111111111111_1111111111111111_1110100001001111_1100101000100000"; -- -0.09253250807523727
	pesos_i(2453) := b"1111111111111111_1111111111111111_1111111100111001_1110111101000110"; -- -0.003022237215191126
	pesos_i(2454) := b"0000000000000000_0000000000000000_0100011001111000_0001111110000000"; -- 0.2752704322338104
	pesos_i(2455) := b"0000000000000000_0000000000000000_0011001101001011_0001101101000000"; -- 0.20036478340625763
	pesos_i(2456) := b"1111111111111111_1111111111111111_1110000000101101_1001101010000000"; -- -0.1243041455745697
	pesos_i(2457) := b"0000000000000000_0000000000000000_0000010001111100_1100110010100000"; -- 0.017529286444187164
	pesos_i(2458) := b"1111111111111111_1111111111111111_1110110100010110_1011101100000000"; -- -0.073871910572052
	pesos_i(2459) := b"1111111111111111_1111111111111111_1011111010010100_0111010000000000"; -- -0.25554728507995605
	pesos_i(2460) := b"1111111111111111_1111111111111111_1010100100110001_0101000010000000"; -- -0.3390912711620331
	pesos_i(2461) := b"0000000000000000_0000000000000000_0100000111010011_1001100100000000"; -- 0.25713497400283813
	pesos_i(2462) := b"0000000000000000_0000000000000000_0100111101100010_1111110110000000"; -- 0.31010422110557556
	pesos_i(2463) := b"0000000000000000_0000000000000000_0101111101110101_0100111110000000"; -- 0.37288376688957214
	pesos_i(2464) := b"1111111111111111_1111111111111111_1100100110111111_1100000100000000"; -- -0.21191781759262085
	pesos_i(2465) := b"1111111111111111_1111111111111111_1111011100101010_1001111010110000"; -- -0.034505922347307205
	pesos_i(2466) := b"0000000000000000_0000000000000000_0001000110001110_1101101100000000"; -- 0.06858605146408081
	pesos_i(2467) := b"0000000000000000_0000000000000000_0110001101000000_0100110010000000"; -- 0.3876998722553253
	pesos_i(2468) := b"1111111111111111_1111111111111111_1111101110011110_1111000011011000"; -- -0.017106005921959877
	pesos_i(2469) := b"0000000000000000_0000000000000000_0000101010101100_1000110011010000"; -- 0.041695404797792435
	pesos_i(2470) := b"0000000000000000_0000000000000000_0010011111101100_1101111100000000"; -- 0.1559581160545349
	pesos_i(2471) := b"0000000000000000_0000000000000000_0100110000000101_1001000010000000"; -- 0.29695990681648254
	pesos_i(2472) := b"0000000000000000_0000000000000000_0001001010001011_0000001010000000"; -- 0.07243362069129944
	pesos_i(2473) := b"0000000000000000_0000000000000000_0000100110001111_1100001010000000"; -- 0.037349849939346313
	pesos_i(2474) := b"1111111111111111_1111111111111111_1111011010010011_0111011100000000"; -- -0.03681236505508423
	pesos_i(2475) := b"0000000000000000_0000000000000000_0011000111000101_1100100110000000"; -- 0.19442424178123474
	pesos_i(2476) := b"0000000000000000_0000000000000000_1000100000110010_0100000100000000"; -- 0.5320168137550354
	pesos_i(2477) := b"0000000000000000_0000000000000000_0010101001001110_0010111001000000"; -- 0.16525544226169586
	pesos_i(2478) := b"0000000000000000_0000000000000000_0111101011100001_1101000110000000"; -- 0.48000821471214294
	pesos_i(2479) := b"0000000000000000_0000000000000000_0101001111000110_1001010000000000"; -- 0.32724881172180176
	pesos_i(2480) := b"1111111111111111_1111111111111111_1110100000001111_0101100011000000"; -- -0.09351582825183868
	pesos_i(2481) := b"1111111111111111_1111111111111111_1111110111111110_0110100011011100"; -- -0.007836767472326756
	pesos_i(2482) := b"0000000000000000_0000000000000000_0000100110101010_1010101111110000"; -- 0.03776049241423607
	pesos_i(2483) := b"0000000000000000_0000000000000000_0101011110011101_0111111110000000"; -- 0.34224697947502136
	pesos_i(2484) := b"0000000000000000_0000000000000000_0010100001000101_0110100101000000"; -- 0.1573091298341751
	pesos_i(2485) := b"1111111111111111_1111111111111111_1101110010011001_1000011110000000"; -- -0.13828232884407043
	pesos_i(2486) := b"1111111111111111_1111111111111111_1110011010010111_0110101011100000"; -- -0.09925205260515213
	pesos_i(2487) := b"0000000000000000_0000000000000000_0101101000110101_1011010100000000"; -- 0.35238200426101685
	pesos_i(2488) := b"0000000000000000_0000000000000000_0100011001011010_0001000010000000"; -- 0.2748117744922638
	pesos_i(2489) := b"0000000000000000_0000000000000000_0110110100100010_1101001110000000"; -- 0.426312655210495
	pesos_i(2490) := b"0000000000000000_0000000000000000_0101010100101011_0010100110000000"; -- 0.3326898515224457
	pesos_i(2491) := b"0000000000000000_0000000000000000_0000011100110101_0100000110111000"; -- 0.028156382963061333
	pesos_i(2492) := b"0000000000000000_0000000000000000_0010110101111100_1111001001000000"; -- 0.17768777906894684
	pesos_i(2493) := b"0000000000000000_0000000000000000_0100111010111001_0101010000000000"; -- 0.30751538276672363
	pesos_i(2494) := b"0000000000000000_0000000000000000_0000001111001101_0001100111110000"; -- 0.014848347753286362
	pesos_i(2495) := b"0000000000000000_0000000000000000_0010110100110000_1000101101000000"; -- 0.17652197182178497
	pesos_i(2496) := b"0000000000000000_0000000000000000_0011010100111110_0000000000000000"; -- 0.207977294921875
	pesos_i(2497) := b"1111111111111111_1111111111111111_1100010010000000_0100011111000000"; -- -0.23241759836673737
	pesos_i(2498) := b"0000000000000000_0000000000000000_0100100001110011_1001010110000000"; -- 0.2830136716365814
	pesos_i(2499) := b"0000000000000000_0000000000000000_0000000110001100_1001101111111010"; -- 0.006051777396351099
	pesos_i(2500) := b"1111111111111111_1111111111111111_1111111011001101_1011011011011100"; -- -0.004673548974096775
	pesos_i(2501) := b"0000000000000000_0000000000000000_0000000001100101_0100011001100001"; -- 0.0015453326050192118
	pesos_i(2502) := b"0000000000000000_0000000000000000_0000100001111011_1010011010110000"; -- 0.0331367664039135
	pesos_i(2503) := b"0000000000000000_0000000000000000_0011010101011101_1111110001000000"; -- 0.2084653526544571
	pesos_i(2504) := b"1111111111111111_1111111111111111_1011110100110011_0100100000000000"; -- -0.26093626022338867
	pesos_i(2505) := b"0000000000000000_0000000000000000_0101000111011010_0001100100000000"; -- 0.3197341561317444
	pesos_i(2506) := b"1111111111111111_1111111111111111_1011000000111101_0101000010000000"; -- -0.3115644156932831
	pesos_i(2507) := b"1111111111111111_1111111111111111_1000000000101001_0011100110000000"; -- -0.4993709623813629
	pesos_i(2508) := b"0000000000000000_0000000000000000_0101111110101111_1101001100000000"; -- 0.3737766146659851
	pesos_i(2509) := b"1111111111111111_1111111111111111_1110110100011111_1101001111000000"; -- -0.07373310625553131
	pesos_i(2510) := b"0000000000000000_0000000000000000_1001111111101100_0110011000000000"; -- 0.6247009038925171
	pesos_i(2511) := b"0000000000000000_0000000000000000_0011011000001110_0111000100000000"; -- 0.21115785837173462
	pesos_i(2512) := b"0000000000000000_0000000000000000_0001110011111000_1111011010000000"; -- 0.11317387223243713
	pesos_i(2513) := b"0000000000000000_0000000000000000_0100110010001100_0110110010000000"; -- 0.29901769757270813
	pesos_i(2514) := b"1111111111111111_1111111111111111_1100011001010000_1110110011000000"; -- -0.22532768547534943
	pesos_i(2515) := b"1111111111111111_1111111111111111_1111111110110111_0100001110000000"; -- -0.001109868404455483
	pesos_i(2516) := b"0000000000000000_0000000000000000_0001111110110110_0001110101100000"; -- 0.12387260049581528
	pesos_i(2517) := b"0000000000000000_0000000000000000_0001000010110010_0100111100100000"; -- 0.06522078067064285
	pesos_i(2518) := b"1111111111111111_1111111111111111_1101110111111010_1101100001000000"; -- -0.13289116322994232
	pesos_i(2519) := b"0000000000000000_0000000000000000_0111010001110001_0000111000000000"; -- 0.45485007762908936
	pesos_i(2520) := b"0000000000000000_0000000000000000_0100100001000110_0110111010000000"; -- 0.2823247015476227
	pesos_i(2521) := b"1111111111111111_1111111111111111_1011100110010100_0111010100000000"; -- -0.2750784754753113
	pesos_i(2522) := b"1111111111111111_1111111111111111_1100100110011000_0001111111000000"; -- -0.21252252161502838
	pesos_i(2523) := b"0000000000000000_0000000000000000_0011011100001101_1010111100000000"; -- 0.2150525450706482
	pesos_i(2524) := b"1111111111111111_1111111111111111_1100101111001100_0101110010000000"; -- -0.20391294360160828
	pesos_i(2525) := b"0000000000000000_0000000000000000_0001101000000001_0000101101000000"; -- 0.10157842934131622
	pesos_i(2526) := b"0000000000000000_0000000000000000_0001000011110111_0111011101100000"; -- 0.06627603620290756
	pesos_i(2527) := b"1111111111111111_1111111111111111_1010101111100010_0101011010000000"; -- -0.32857760787010193
	pesos_i(2528) := b"0000000000000000_0000000000000000_0100111110001000_0011000110000000"; -- 0.3106718957424164
	pesos_i(2529) := b"1111111111111111_1111111111111111_1101000110110001_0111010011000000"; -- -0.18088598549365997
	pesos_i(2530) := b"0000000000000000_0000000000000000_0010100111101010_1111111110000000"; -- 0.1637420356273651
	pesos_i(2531) := b"0000000000000000_0000000000000000_0000000000111110_0000101100000110"; -- 0.000946702086366713
	pesos_i(2532) := b"0000000000000000_0000000000000000_0011010000011000_1110110000000000"; -- 0.203505277633667
	pesos_i(2533) := b"0000000000000000_0000000000000000_0011011110010001_0011100010000000"; -- 0.2170596420764923
	pesos_i(2534) := b"0000000000000000_0000000000000000_0011101110100111_1001110000000000"; -- 0.23302626609802246
	pesos_i(2535) := b"1111111111111111_1111111111111111_1100111100100110_0100101011000000"; -- -0.19082196056842804
	pesos_i(2536) := b"1111111111111111_1111111111111111_1111101011010111_1011001000111000"; -- -0.020146237686276436
	pesos_i(2537) := b"1111111111111111_1111111111111111_1110101011101011_0100111011000000"; -- -0.08234699070453644
	pesos_i(2538) := b"0000000000000000_0000000000000000_1000100100101001_0100011100000000"; -- 0.5357860922813416
	pesos_i(2539) := b"0000000000000000_0000000000000000_0000000001100101_1010110111101111"; -- 0.0015515049453824759
	pesos_i(2540) := b"1111111111111111_1111111111111111_1100000011100100_0101111011000000"; -- -0.24651534855365753
	pesos_i(2541) := b"0000000000000000_0000000000000000_0001000110010011_0110110010100000"; -- 0.06865576654672623
	pesos_i(2542) := b"1111111111111111_1111111111111111_1100100001101100_1111010000000000"; -- -0.2170875072479248
	pesos_i(2543) := b"0000000000000000_0000000000000000_1000101011000101_1010100000000000"; -- 0.5420784950256348
	pesos_i(2544) := b"1111111111111111_1111111111111111_1100110011001101_1101111101000000"; -- -0.1999836415052414
	pesos_i(2545) := b"1111111111111111_1111111111111111_1110010111100111_1000000010000000"; -- -0.10193631052970886
	pesos_i(2546) := b"1111111111111111_1111111111111111_1001111100000001_0010010010000000"; -- -0.3788888156414032
	pesos_i(2547) := b"0000000000000000_0000000000000000_0011001101010011_0110000100000000"; -- 0.2004910111427307
	pesos_i(2548) := b"0000000000000000_0000000000000000_0100100001101000_0011000000000000"; -- 0.2828397750854492
	pesos_i(2549) := b"0000000000000000_0000000000000000_0010001011000111_0101100000000000"; -- 0.13585424423217773
	pesos_i(2550) := b"1111111111111111_1111111111111111_1110011100010111_1100100001000000"; -- -0.09729336202144623
	pesos_i(2551) := b"1111111111111111_1111111111111111_1100010010011010_0101011111000000"; -- -0.23201991617679596
	pesos_i(2552) := b"1111111111111111_1111111111111111_1001100010111001_0111110110000000"; -- -0.4034196436405182
	pesos_i(2553) := b"1111111111111111_1111111111111111_1110011110011000_0010110100000000"; -- -0.09533423185348511
	pesos_i(2554) := b"0000000000000000_0000000000000000_0000000001000100_0000010111110111"; -- 0.0010379531886428595
	pesos_i(2555) := b"1111111111111111_1111111111111111_1110011110110111_1010111000100000"; -- -0.09485351294279099
	pesos_i(2556) := b"0000000000000000_0000000000000000_0100100010011010_0110000100000000"; -- 0.2836056351661682
	pesos_i(2557) := b"0000000000000000_0000000000000000_0000000000001110_0001011110011000"; -- 0.000215029256651178
	pesos_i(2558) := b"0000000000000000_0000000000000000_0000000000001001_0000010101101101"; -- 0.00013765260518994182
	pesos_i(2559) := b"0000000000000000_0000000000000000_0001000100010010_0100101100100000"; -- 0.06668538600206375
	pesos_i(2560) := b"1111111111111111_1111111111111111_1000010010100111_0011101100000000"; -- -0.48182326555252075
	pesos_i(2561) := b"0000000000000000_0000000000000000_0101011001010100_1110001110000000"; -- 0.3372327983379364
	pesos_i(2562) := b"0000000000000000_0000000000000000_1000010011111001_1110000100000000"; -- 0.519437849521637
	pesos_i(2563) := b"1111111111111111_1111111111111111_1010000100001011_1001101110000000"; -- -0.3709166347980499
	pesos_i(2564) := b"1111111111111111_1111111111111111_1011011011000001_0101000000000000"; -- -0.28611278533935547
	pesos_i(2565) := b"0000000000000000_0000000000000000_0101001010000000_1001111110000000"; -- 0.3222751319408417
	pesos_i(2566) := b"1111111111111111_1111111111111111_1111101111000000_0111101100011000"; -- -0.01659422554075718
	pesos_i(2567) := b"0000000000000000_0000000000000000_0111000111100111_1110000110000000"; -- 0.44494447112083435
	pesos_i(2568) := b"0000000000000000_0000000000000000_0000101001101010_0001011000000000"; -- 0.04068124294281006
	pesos_i(2569) := b"1111111111111111_1111111111111111_1110011000101100_0011100000100000"; -- -0.10088776797056198
	pesos_i(2570) := b"1111111111111111_1111111111111111_1111010111001111_1101001011010000"; -- -0.03979761525988579
	pesos_i(2571) := b"0000000000000000_0000000000000000_0111010100101110_1110100000000000"; -- 0.4577469825744629
	pesos_i(2572) := b"1111111111111111_1111111111111111_1101100010000011_1001011100000000"; -- -0.15424209833145142
	pesos_i(2573) := b"1111111111111111_1111111111111111_1010010100001000_0000011010000000"; -- -0.35534629225730896
	pesos_i(2574) := b"0000000000000000_0000000000000000_0001101100111111_0010001100000000"; -- 0.10643213987350464
	pesos_i(2575) := b"0000000000000000_0000000000000000_0110010011000111_1001011000000000"; -- 0.3936704397201538
	pesos_i(2576) := b"1111111111111111_1111111111111111_1010110100000000_0000101000000000"; -- -0.32421815395355225
	pesos_i(2577) := b"1111111111111111_1111111111111111_1110011100001010_1101011110100000"; -- -0.0974908098578453
	pesos_i(2578) := b"0000000000000000_0000000000000000_0100010000101010_1110100000000000"; -- 0.2662796974182129
	pesos_i(2579) := b"0000000000000000_0000000000000000_0110000111100011_1010101010000000"; -- 0.3823801577091217
	pesos_i(2580) := b"1111111111111111_1111111111111111_1001111001111010_0110000000000000"; -- -0.38094520568847656
	pesos_i(2581) := b"0000000000000000_0000000000000000_0000111010101000_1000010000100000"; -- 0.05725885182619095
	pesos_i(2582) := b"0000000000000000_0000000000000000_1001001001100001_0101111000000000"; -- 0.5717982053756714
	pesos_i(2583) := b"0000000000000000_0000000000000000_0000011100010110_1011001101000000"; -- 0.02769012749195099
	pesos_i(2584) := b"1111111111111111_1111111111111111_1101100011011110_1000010100000000"; -- -0.15285462141036987
	pesos_i(2585) := b"0000000000000000_0000000000000000_0001111101011010_0100001101000000"; -- 0.12247104942798615
	pesos_i(2586) := b"0000000000000000_0000000000000000_0110100101100000_1100010000000000"; -- 0.411632776260376
	pesos_i(2587) := b"0000000000000000_0000000000000000_0101100110110111_1101110010000000"; -- 0.3504617512226105
	pesos_i(2588) := b"1111111111111111_1111111111111111_0111111100001111_0001100000000000"; -- -0.5036759376525879
	pesos_i(2589) := b"1111111111111111_1111111111111111_1100010011011110_0101010001000000"; -- -0.23098252713680267
	pesos_i(2590) := b"0000000000000000_0000000000000000_0111100000000111_0110110100000000"; -- 0.468863308429718
	pesos_i(2591) := b"0000000000000000_0000000000000000_0001011101101110_1110011001100000"; -- 0.09153594821691513
	pesos_i(2592) := b"1111111111111111_1111111111111110_1110000110010110_0000011000000000"; -- -1.1188045740127563
	pesos_i(2593) := b"1111111111111111_1111111111111111_1110111010000110_0001110010000000"; -- -0.0682661235332489
	pesos_i(2594) := b"0000000000000000_0000000000000000_0011111101000101_0001011011000000"; -- 0.24714796245098114
	pesos_i(2595) := b"1111111111111111_1111111111111111_1111110111100110_0010111011110000"; -- -0.008206430822610855
	pesos_i(2596) := b"0000000000000000_0000000000000000_0111011101101111_1100100000000000"; -- 0.4665493965148926
	pesos_i(2597) := b"1111111111111111_1111111111111111_1110010101000110_1011100010100000"; -- -0.10438963025808334
	pesos_i(2598) := b"1111111111111111_1111111111111111_1011110110100101_0000010110000000"; -- -0.25920072197914124
	pesos_i(2599) := b"0000000000000000_0000000000000000_0000010111101000_0000011110100000"; -- 0.023071743547916412
	pesos_i(2600) := b"1111111111111111_1111111111111111_1101001110010111_1000100000000000"; -- -0.17346906661987305
	pesos_i(2601) := b"0000000000000000_0000000000000000_0011101101000010_1111011010000000"; -- 0.23149052262306213
	pesos_i(2602) := b"0000000000000000_0000000000000000_0110001010001010_1100000100000000"; -- 0.38492971658706665
	pesos_i(2603) := b"0000000000000000_0000000000000000_0111101001100111_0100110010000000"; -- 0.4781387150287628
	pesos_i(2604) := b"0000000000000000_0000000000000000_1100011011100011_1001011000000000"; -- 0.7769101858139038
	pesos_i(2605) := b"0000000000000000_0000000000000000_0111110101011001_1111010000000000"; -- 0.4896538257598877
	pesos_i(2606) := b"0000000000000000_0000000000000000_0010011011111111_0110101011000000"; -- 0.15233485400676727
	pesos_i(2607) := b"0000000000000000_0000000000000000_0011000110010110_0011110101000000"; -- 0.1936987191438675
	pesos_i(2608) := b"0000000000000000_0000000000000000_0110000000000010_1110011110000000"; -- 0.3750443160533905
	pesos_i(2609) := b"0000000000000000_0000000000000000_0111010101110001_0100110100000000"; -- 0.4587600827217102
	pesos_i(2610) := b"1111111111111111_1111111111111111_1100111100000011_0001100110000000"; -- -0.19135895371437073
	pesos_i(2611) := b"1111111111111111_1111111111111111_0001100101110000_1100011000000000"; -- -0.9006229639053345
	pesos_i(2612) := b"0000000000000000_0000000000000000_0011110001011000_0000101011000000"; -- 0.23571841418743134
	pesos_i(2613) := b"0000000000000000_0000000000000000_0000110111000111_0110100101110000"; -- 0.053824033588171005
	pesos_i(2614) := b"1111111111111111_1111111111111111_1010111100000100_1010011000000000"; -- -0.3163353204727173
	pesos_i(2615) := b"0000000000000000_0000000000000000_0011101111000110_0011101011000000"; -- 0.23349349200725555
	pesos_i(2616) := b"1111111111111111_1111111111111111_1010110011110011_1001111100000000"; -- -0.3244076371192932
	pesos_i(2617) := b"0000000000000000_0000000000000000_0111101010100100_1101110000000000"; -- 0.4790780544281006
	pesos_i(2618) := b"0000000000000000_0000000000000000_0010000101100110_1111011111000000"; -- 0.1304774135351181
	pesos_i(2619) := b"0000000000000000_0000000000000000_0011010000010110_0111010001000000"; -- 0.20346762239933014
	pesos_i(2620) := b"0000000000000000_0000000000000000_0001011001101011_1001001100000000"; -- 0.08757895231246948
	pesos_i(2621) := b"1111111111111111_1111111111111111_1001111010001110_0011111100000000"; -- -0.38064199686050415
	pesos_i(2622) := b"1111111111111111_1111111111111111_1110010111010101_0011110000000000"; -- -0.10221505165100098
	pesos_i(2623) := b"1111111111111111_1111111111111111_0100001010110110_0000110000000000"; -- -0.7394096851348877
	pesos_i(2624) := b"1111111111111111_1111111111111111_1101101000110101_0001111111000000"; -- -0.14762689173221588
	pesos_i(2625) := b"0000000000000000_0000000000000000_0100101100110010_1011001010000000"; -- 0.2937423288822174
	pesos_i(2626) := b"0000000000000000_0000000000000000_0001111010110011_1100001110100000"; -- 0.11993048340082169
	pesos_i(2627) := b"0000000000000000_0000000000000000_0000111110011011_0100100010100000"; -- 0.06096319109201431
	pesos_i(2628) := b"1111111111111111_1111111111111111_1111100111001101_1001100101000000"; -- -0.02420656383037567
	pesos_i(2629) := b"0000000000000000_0000000000000000_0011000001101110_1010001000000000"; -- 0.1891881227493286
	pesos_i(2630) := b"0000000000000000_0000000000000000_1100001111101100_0001101000000000"; -- 0.7653213739395142
	pesos_i(2631) := b"1111111111111111_1111111111111111_1001101110111000_0010011000000000"; -- -0.39172136783599854
	pesos_i(2632) := b"1111111111111111_1111111111111111_1111101100101101_1001101010100000"; -- -0.018835388123989105
	pesos_i(2633) := b"0000000000000000_0000000000000000_1011110100100100_1001111000000000"; -- 0.7388399839401245
	pesos_i(2634) := b"0000000000000000_0000000000000000_0011000100101111_0110001110000000"; -- 0.19212934374809265
	pesos_i(2635) := b"1111111111111111_1111111111111111_1001101010101101_1100111010000000"; -- -0.3957854211330414
	pesos_i(2636) := b"0000000000000000_0000000000000000_0001111111000101_0111110101000000"; -- 0.12410719692707062
	pesos_i(2637) := b"0000000000000000_0000000000000000_0100100011110100_0100011110000000"; -- 0.28497740626335144
	pesos_i(2638) := b"1111111111111111_1111111111111111_1100000001111111_1110111100000000"; -- -0.24804788827896118
	pesos_i(2639) := b"0000000000000000_0000000000000000_1000011111111001_0101000000000000"; -- 0.5311479568481445
	pesos_i(2640) := b"1111111111111111_1111111111111111_1100110010000011_0011100101000000"; -- -0.2011226862668991
	pesos_i(2641) := b"1111111111111111_1111111111111111_1110100100100111_1101000101100000"; -- -0.08923617750406265
	pesos_i(2642) := b"1111111111111111_1111111111111111_1100001111101001_0110101010000000"; -- -0.23471960425376892
	pesos_i(2643) := b"1111111111111111_1111111111111111_1001000110000111_1111101010000000"; -- -0.43151888251304626
	pesos_i(2644) := b"1111111111111111_1111111111111111_1011000111110010_1101000010000000"; -- -0.30488869547843933
	pesos_i(2645) := b"1111111111111111_1111111111111111_1111111110100101_0001110101100000"; -- -0.001386798918247223
	pesos_i(2646) := b"0000000000000000_0000000000000000_0001011110000110_0001011000000000"; -- 0.09188973903656006
	pesos_i(2647) := b"0000000000000000_0000000000000000_0011011011010101_1001111111000000"; -- 0.21419714391231537
	pesos_i(2648) := b"0000000000000000_0000000000000000_0111010100101010_0011011010000000"; -- 0.45767536759376526
	pesos_i(2649) := b"1111111111111111_1111111111111111_1011001010000001_0010000100000000"; -- -0.3027171492576599
	pesos_i(2650) := b"0000000000000000_0000000000000000_0000000110110101_0110101011110110"; -- 0.00667446618899703
	pesos_i(2651) := b"0000000000000000_0000000000000000_0110110111001101_0001101010000000"; -- 0.42891088128089905
	pesos_i(2652) := b"0000000000000000_0000000000000000_0001110001001111_0010111010100000"; -- 0.11058322340250015
	pesos_i(2653) := b"1111111111111111_1111111111111111_1111000110010010_0101100010100000"; -- -0.05636068433523178
	pesos_i(2654) := b"0000000000000000_0000000000000000_0000010101011001_1101000001001000"; -- 0.020901696756482124
	pesos_i(2655) := b"0000000000000000_0000000000000000_0011101011010000_0110111000000000"; -- 0.2297428846359253
	pesos_i(2656) := b"0000000000000000_0000000000000000_0101001101110010_1000100100000000"; -- 0.32596641778945923
	pesos_i(2657) := b"1111111111111111_1111111111111111_1110101111100101_0001100111100000"; -- -0.07853544503450394
	pesos_i(2658) := b"0000000000000000_0000000000000000_0100001110100011_1110001110000000"; -- 0.2642194926738739
	pesos_i(2659) := b"1111111111111111_1111111111111111_1101100010111011_0000101111000000"; -- -0.1533959060907364
	pesos_i(2660) := b"0000000000000000_0000000000000000_0110001000111010_0001001100000000"; -- 0.38369864225387573
	pesos_i(2661) := b"0000000000000000_0000000000000000_0001000110011100_1100010011000000"; -- 0.06879834830760956
	pesos_i(2662) := b"1111111111111111_1111111111111111_1111010111101111_0101000110000000"; -- -0.039317041635513306
	pesos_i(2663) := b"0000000000000000_0000000000000000_0001111011110111_1101010110000000"; -- 0.12096914649009705
	pesos_i(2664) := b"1111111111111111_1111111111111111_0111100110001001_0001011000000000"; -- -0.5252519845962524
	pesos_i(2665) := b"0000000000000000_0000000000000000_0110001111001000_0010101010000000"; -- 0.38977304100990295
	pesos_i(2666) := b"0000000000000000_0000000000000000_0000010111000110_0001000110010000"; -- 0.022553537040948868
	pesos_i(2667) := b"1111111111111111_1111111111111111_1110111000111001_0010001110100000"; -- -0.06944062560796738
	pesos_i(2668) := b"0000000000000000_0000000000000000_0010110011010110_0001101110000000"; -- 0.17514201998710632
	pesos_i(2669) := b"1111111111111111_1111111111111111_1101101001110010_1000110111000000"; -- -0.1466895490884781
	pesos_i(2670) := b"0000000000000000_0000000000000000_0110000000100010_1101111000000000"; -- 0.37553203105926514
	pesos_i(2671) := b"0000000000000000_0000000000000000_1000000100011010_1011111100000000"; -- 0.5043143630027771
	pesos_i(2672) := b"1111111111111111_1111111111111111_1101111101000111_0111100101000000"; -- -0.12781564891338348
	pesos_i(2673) := b"0000000000000000_0000000000000000_0100100101000101_0000110000000000"; -- 0.2862098217010498
	pesos_i(2674) := b"1111111111111111_1111111111111111_1000010000000010_1000110110000000"; -- -0.4843360483646393
	pesos_i(2675) := b"1111111111111111_1111111111111111_1100001101111001_1001011101000000"; -- -0.23642592132091522
	pesos_i(2676) := b"1111111111111111_1111111111111111_1110001010110000_0001010000000000"; -- -0.11450076103210449
	pesos_i(2677) := b"1111111111111111_1111111111111111_1101111100000010_0100010111000000"; -- -0.12887157499790192
	pesos_i(2678) := b"0000000000000000_0000000000000000_0000100101011011_1011000100100000"; -- 0.03655535727739334
	pesos_i(2679) := b"0000000000000000_0000000000000000_0110011110111001_0101000110000000"; -- 0.4051714837551117
	pesos_i(2680) := b"1111111111111111_1111111111111111_1101011100101001_0100001001000000"; -- -0.15952669084072113
	pesos_i(2681) := b"0000000000000000_0000000000000000_0100111001100110_0010001110000000"; -- 0.3062460124492645
	pesos_i(2682) := b"1111111111111111_1111111111111111_1110001001111111_1001111110100000"; -- -0.11524011939764023
	pesos_i(2683) := b"0000000000000000_0000000000000000_0010010011010100_0001011101000000"; -- 0.14386124908924103
	pesos_i(2684) := b"0000000000000000_0000000000000000_0010000101001010_1010111000000000"; -- 0.13004577159881592
	pesos_i(2685) := b"0000000000000000_0000000000000000_0011010011101000_1001000011000000"; -- 0.20667366683483124
	pesos_i(2686) := b"1111111111111111_1111111111111111_1110110101110001_1000100111000000"; -- -0.07248629629611969
	pesos_i(2687) := b"0000000000000000_0000000000000000_1000000000111010_0001001100000000"; -- 0.5008861422538757
	pesos_i(2688) := b"1111111111111111_1111111111111111_1101000110111010_1100000001000000"; -- -0.18074415624141693
	pesos_i(2689) := b"0000000000000000_0000000000000000_0100011101110011_0110111110000000"; -- 0.27910515666007996
	pesos_i(2690) := b"0000000000000000_0000000000000000_0100010001001010_0100010000000000"; -- 0.2667582035064697
	pesos_i(2691) := b"1111111111111111_1111111111111111_1111011100101110_0100000111110000"; -- -0.03445041552186012
	pesos_i(2692) := b"0000000000000000_0000000000000000_0110000001011101_0001100100000000"; -- 0.3764205574989319
	pesos_i(2693) := b"0000000000000000_0000000000000000_1001001110010110_0011001000000000"; -- 0.5765105485916138
	pesos_i(2694) := b"1111111111111111_1111111111111111_1110100011010010_1101101110000000"; -- -0.0905325710773468
	pesos_i(2695) := b"1111111111111111_1111111111111111_1111110000000101_1110111001011000"; -- -0.015534499660134315
	pesos_i(2696) := b"0000000000000000_0000000000000000_0010110110110100_1111001001000000"; -- 0.17854227125644684
	pesos_i(2697) := b"0000000000000000_0000000000000000_0001110001010101_1001001011000000"; -- 0.11068074405193329
	pesos_i(2698) := b"0000000000000000_0000000000000000_0011100001100100_0001111101000000"; -- 0.22027774155139923
	pesos_i(2699) := b"1111111111111111_1111111111111111_1101110011011001_1111001001000000"; -- -0.13729940354824066
	pesos_i(2700) := b"1111111111111111_1111111111111111_1011001100111111_0110010000000000"; -- -0.29981398582458496
	pesos_i(2701) := b"0000000000000000_0000000000000000_0000110110110111_0111100111000000"; -- 0.053580865263938904
	pesos_i(2702) := b"0000000000000000_0000000000000000_0000111001110100_0100110011110000"; -- 0.05646210536360741
	pesos_i(2703) := b"0000000000000000_0000000000000000_0010101010111000_0010100010000000"; -- 0.1668725311756134
	pesos_i(2704) := b"1111111111111111_1111111111111111_1110100110110110_0010001010100000"; -- -0.08706458657979965
	pesos_i(2705) := b"1111111111111111_1111111111111111_1100111010000010_1010101101000000"; -- -0.19331865012645721
	pesos_i(2706) := b"0000000000000000_0000000000000000_0011001111000010_1011010010000000"; -- 0.20218971371650696
	pesos_i(2707) := b"0000000000000000_0000000000000000_0010011101010011_1101001001000000"; -- 0.15362276136875153
	pesos_i(2708) := b"1111111111111111_1111111111111111_1110101101010110_0100000101100000"; -- -0.08071509748697281
	pesos_i(2709) := b"0000000000000000_0000000000000000_0011011001010010_0011001001000000"; -- 0.21219171583652496
	pesos_i(2710) := b"0000000000000000_0000000000000000_0001110010000000_0100100011100000"; -- 0.111332468688488
	pesos_i(2711) := b"1111111111111111_1111111111111111_1110111001010011_0110000010000000"; -- -0.06904026865959167
	pesos_i(2712) := b"0000000000000000_0000000000000000_0110101010101110_0100111100000000"; -- 0.41672223806381226
	pesos_i(2713) := b"0000000000000000_0000000000000000_0110101110010111_1111110010000000"; -- 0.4202878773212433
	pesos_i(2714) := b"1111111111111111_1111111111111111_1111010001111101_0001110101110000"; -- -0.044965896755456924
	pesos_i(2715) := b"0000000000000000_0000000000000000_0000101100110000_0111001001100000"; -- 0.043707989156246185
	pesos_i(2716) := b"1111111111111111_1111111111111111_1100011001101000_1001111111000000"; -- -0.22496606409549713
	pesos_i(2717) := b"0000000000000000_0000000000000000_0001001101110011_1100001111100000"; -- 0.07598518580198288
	pesos_i(2718) := b"0000000000000000_0000000000000000_0011111110001101_0101001111000000"; -- 0.24825023114681244
	pesos_i(2719) := b"0000000000000000_0000000000000000_0000010111100001_0100101111101000"; -- 0.022969001904129982
	pesos_i(2720) := b"1111111111111111_1111111111111111_1011011000000101_0001011100000000"; -- -0.28898483514785767
	pesos_i(2721) := b"0000000000000000_0000000000000000_0010010010110111_0101101100000000"; -- 0.14342278242111206
	pesos_i(2722) := b"0000000000000000_0000000000000000_0000000010010011_1000010110101110"; -- 0.0022510099224746227
	pesos_i(2723) := b"0000000000000000_0000000000000000_0001000000000001_0111100101100000"; -- 0.06252249330282211
	pesos_i(2724) := b"1111111111111111_1111111111111111_1111010100100001_1011111011110000"; -- -0.0424538291990757
	pesos_i(2725) := b"1111111111111111_1111111111111111_1011110110111010_1010001010000000"; -- -0.258870929479599
	pesos_i(2726) := b"1111111111111111_1111111111111111_1110111011101111_0001000110100000"; -- -0.06666459888219833
	pesos_i(2727) := b"0000000000000000_0000000000000000_0001000100001001_0110100110000000"; -- 0.0665498673915863
	pesos_i(2728) := b"1111111111111111_1111111111111111_1111001111010001_1000011110010000"; -- -0.047584082931280136
	pesos_i(2729) := b"1111111111111111_1111111111111111_1110101100110000_0000010010100000"; -- -0.08129855245351791
	pesos_i(2730) := b"1111111111111111_1111111111111111_1101000001001001_0001011110000000"; -- -0.18638470768928528
	pesos_i(2731) := b"1111111111111111_1111111111111111_1001010110101000_1100100010000000"; -- -0.41539332270622253
	pesos_i(2732) := b"1111111111111111_1111111111111111_1111001101101100_1010010110010000"; -- -0.049123432487249374
	pesos_i(2733) := b"0000000000000000_0000000000000000_0100000000010110_0001110010000000"; -- 0.2503373920917511
	pesos_i(2734) := b"1111111111111111_1111111111111111_1111111011011000_1101101011010110"; -- -0.004503557924181223
	pesos_i(2735) := b"0000000000000000_0000000000000000_0001100110001001_0000001001100000"; -- 0.09974684566259384
	pesos_i(2736) := b"0000000000000000_0000000000000000_0010011011100111_0101000010000000"; -- 0.15196707844734192
	pesos_i(2737) := b"0000000000000000_0000000000000000_0000110111011100_1111110010100000"; -- 0.05415324121713638
	pesos_i(2738) := b"0000000000000000_0000000000000000_0001111110011000_0001000100100000"; -- 0.12341410666704178
	pesos_i(2739) := b"1111111111111111_1111111111111110_1011110010100011_1110001000000000"; -- -1.2631243467330933
	pesos_i(2740) := b"0000000000000000_0000000000000000_0011111011110101_1101001010000000"; -- 0.24593845009803772
	pesos_i(2741) := b"0000000000000000_0000000000000000_0000110111000101_1010101111110000"; -- 0.05379747971892357
	pesos_i(2742) := b"0000000000000000_0000000000000000_0000110000101110_0000011010010000"; -- 0.04757729545235634
	pesos_i(2743) := b"0000000000000000_0000000000000000_0111001110011010_1000000000000000"; -- 0.45157623291015625
	pesos_i(2744) := b"0000000000000000_0000000000000000_0010000000011011_0111111011000000"; -- 0.12541954219341278
	pesos_i(2745) := b"1111111111111111_1111111111111111_1110100100101011_1000001011000000"; -- -0.08917982876300812
	pesos_i(2746) := b"0000000000000000_0000000000000000_0001101110001011_0101001110000000"; -- 0.10759469866752625
	pesos_i(2747) := b"0000000000000000_0000000000000000_0000110110111101_0000000011110000"; -- 0.05366521701216698
	pesos_i(2748) := b"0000000000000000_0000000000000000_0100000000010011_1001111000000000"; -- 0.250299334526062
	pesos_i(2749) := b"1111111111111111_1111111111111111_1110110100010110_0010001011100000"; -- -0.07388097792863846
	pesos_i(2750) := b"0000000000000000_0000000000000000_0100100100010110_1000110000000000"; -- 0.28550028800964355
	pesos_i(2751) := b"1111111111111111_1111111111111111_0010001001110110_0011001000000000"; -- -0.8653839826583862
	pesos_i(2752) := b"0000000000000000_0000000000000000_0010000110001110_0111110100000000"; -- 0.13108044862747192
	pesos_i(2753) := b"0000000000000000_0000000000000000_0110010001100110_0010001100000000"; -- 0.39218348264694214
	pesos_i(2754) := b"1111111111111111_1111111111111111_1100100111101001_1001000110000000"; -- -0.21127977967262268
	pesos_i(2755) := b"0000000000000000_0000000000000000_0100011101011110_1010010110000000"; -- 0.2787879407405853
	pesos_i(2756) := b"0000000000000000_0000000000000000_0101011011100110_0010110110000000"; -- 0.3394497334957123
	pesos_i(2757) := b"1111111111111111_1111111111111111_1101001101000001_0011011011000000"; -- -0.17478616535663605
	pesos_i(2758) := b"0000000000000000_0000000000000000_0110111111001011_0110011110000000"; -- 0.43669745326042175
	pesos_i(2759) := b"0000000000000000_0000000000000000_0011110000101101_1101001100000000"; -- 0.2350742220878601
	pesos_i(2760) := b"0000000000000000_0000000000000000_0011011000010011_1100001110000000"; -- 0.2112390697002411
	pesos_i(2761) := b"0000000000000000_0000000000000000_0110010101010111_1111100000000000"; -- 0.3958735466003418
	pesos_i(2762) := b"1111111111111111_1111111111111111_1111011111100010_0111000000100000"; -- -0.03170108050107956
	pesos_i(2763) := b"1111111111111111_1111111111111111_1011111010011111_1101010010000000"; -- -0.25537368655204773
	pesos_i(2764) := b"0000000000000000_0000000000000000_0000011100000110_0100010111010000"; -- 0.027439463883638382
	pesos_i(2765) := b"0000000000000000_0000000000000000_0101011010101101_1001011100000000"; -- 0.3385862708091736
	pesos_i(2766) := b"1111111111111111_1111111111111111_1010001111111011_1000011110000000"; -- -0.35944321751594543
	pesos_i(2767) := b"1111111111111111_1111111111111111_1011101001011011_0011010100000000"; -- -0.2720457911491394
	pesos_i(2768) := b"0000000000000000_0000000000000000_0011010101110010_0001110010000000"; -- 0.2087724506855011
	pesos_i(2769) := b"1111111111111111_1111111111111111_0010110011101101_1011111100000000"; -- -0.8244972825050354
	pesos_i(2770) := b"1111111111111111_1111111111111111_1100111110111000_1011110011000000"; -- -0.18858738243579865
	pesos_i(2771) := b"1111111111111111_1111111111111111_1101100100001111_1001010001000000"; -- -0.15210603177547455
	pesos_i(2772) := b"0000000000000000_0000000000000000_0011110011101110_1100010111000000"; -- 0.23801837861537933
	pesos_i(2773) := b"0000000000000000_0000000000000000_0111000111100011_1011001010000000"; -- 0.4448806345462799
	pesos_i(2774) := b"0000000000000000_0000000000000000_1000000000010001_1011011000000000"; -- 0.5002702474594116
	pesos_i(2775) := b"0000000000000000_0000000000000000_0001111011010111_0010000110000000"; -- 0.12047013640403748
	pesos_i(2776) := b"0000000000000000_0000000000000000_0010011100101000_0100110111000000"; -- 0.1529587358236313
	pesos_i(2777) := b"0000000000000000_0000000000000000_0001100001010110_1111111000000000"; -- 0.09507739543914795
	pesos_i(2778) := b"0000000000000000_0000000000000000_0101010101011100_0000001010000000"; -- 0.33343520760536194
	pesos_i(2779) := b"0000000000000000_0000000000000000_0010111110101000_1100111110000000"; -- 0.1861695945262909
	pesos_i(2780) := b"0000000000000000_0000000000000000_0010101010011101_0011110111000000"; -- 0.16646181046962738
	pesos_i(2781) := b"0000000000000000_0000000000000000_0011000110001101_0101000011000000"; -- 0.1935625523328781
	pesos_i(2782) := b"1111111111111111_1111111111111111_1100001101110110_1111011000000000"; -- -0.23646605014801025
	pesos_i(2783) := b"0000000000000000_0000000000000000_0000110101000011_0010111011010000"; -- 0.05180637910962105
	pesos_i(2784) := b"1111111111111111_1111111111111111_1111111011000000_1001010101010100"; -- -0.0048739118501544
	pesos_i(2785) := b"1111111111111111_1111111111111111_1110110010110000_0101100100100000"; -- -0.0754341408610344
	pesos_i(2786) := b"0000000000000000_0000000000000000_0011001101100111_1010000100000000"; -- 0.20080000162124634
	pesos_i(2787) := b"1111111111111111_1111111111111111_1110010100011111_1101001000100000"; -- -0.10498320311307907
	pesos_i(2788) := b"0000000000000000_0000000000000000_0101111111111110_0000101100000000"; -- 0.37497013807296753
	pesos_i(2789) := b"0000000000000000_0000000000000000_0010010100111100_1010111101000000"; -- 0.1454572230577469
	pesos_i(2790) := b"0000000000000000_0000000000000000_0000110100000110_0111000010110000"; -- 0.05087951943278313
	pesos_i(2791) := b"0000000000000000_0000000000000000_0110010011010111_0111011010000000"; -- 0.3939127027988434
	pesos_i(2792) := b"1111111111111111_1111111111111111_1111011001111100_0011110000000000"; -- -0.03716683387756348
	pesos_i(2793) := b"0000000000000000_0000000000000000_0010000110101011_0000101001000000"; -- 0.13151611387729645
	pesos_i(2794) := b"1111111111111111_1111111111111111_1100000100101000_1000100011000000"; -- -0.24547524750232697
	pesos_i(2795) := b"0000000000000000_0000000000000000_0001001110111010_1111100000100000"; -- 0.0770716741681099
	pesos_i(2796) := b"1111111111111111_1111111111111111_0110101100010000_0010011000000000"; -- -0.5817848443984985
	pesos_i(2797) := b"1111111111111111_1111111111111111_1110111001010011_0100100010000000"; -- -0.06904169917106628
	pesos_i(2798) := b"0000000000000000_0000000000000000_0011101011001100_1011100010000000"; -- 0.22968629002571106
	pesos_i(2799) := b"0000000000000000_0000000000000000_0011111001000000_0110000011000000"; -- 0.24316982924938202
	pesos_i(2800) := b"0000000000000000_0000000000000000_0010001011111100_1001100001000000"; -- 0.13666678965091705
	pesos_i(2801) := b"0000000000000000_0000000000000000_0100001101000001_0000000000000000"; -- 0.2627105712890625
	pesos_i(2802) := b"1111111111111111_1111111111111111_1101001101100000_0110011101000000"; -- -0.17431025207042694
	pesos_i(2803) := b"0000000000000000_0000000000000000_0100000000110011_1100111010000000"; -- 0.2507905066013336
	pesos_i(2804) := b"1111111111111111_1111111111111111_1111010110110000_1101011001010000"; -- -0.040270429104566574
	pesos_i(2805) := b"1111111111111111_1111111111111111_1010001110100010_0111100010000000"; -- -0.36080214381217957
	pesos_i(2806) := b"0000000000000000_0000000000000000_0011010100100100_0011011110000000"; -- 0.20758387446403503
	pesos_i(2807) := b"1111111111111111_1111111111111111_1111011000011110_1011010101010000"; -- -0.03859392926096916
	pesos_i(2808) := b"1111111111111111_1111111111111111_1110000100000001_0011110110000000"; -- -0.12107482552528381
	pesos_i(2809) := b"1111111111111111_1111111111111111_1111101001110010_1001100000010000"; -- -0.021688934415578842
	pesos_i(2810) := b"1111111111111111_1111111111111111_1101111011001101_1111000011000000"; -- -0.12967009842395782
	pesos_i(2811) := b"0000000000000000_0000000000000000_0011101000011110_1001000010000000"; -- 0.22702887654304504
	pesos_i(2812) := b"1111111111111111_1111111111111111_1001011100110101_0110010110000000"; -- -0.4093414843082428
	pesos_i(2813) := b"0000000000000000_0000000000000000_0000001011100101_1001101111000000"; -- 0.011316046118736267
	pesos_i(2814) := b"0000000000000000_0000000000000000_0001101101001001_0010111101100000"; -- 0.10658546537160873
	pesos_i(2815) := b"0000000000000000_0000000000000000_0101001110101101_0100001100000000"; -- 0.32686251401901245
	pesos_i(2816) := b"1111111111111111_1111111111111111_1111010001011000_0000110000000000"; -- -0.045531511306762695
	pesos_i(2817) := b"0000000000000000_0000000000000000_0100001110101000_0101000000000000"; -- 0.26428699493408203
	pesos_i(2818) := b"1111111111111111_1111111111111111_1111100101101111_1101000001100000"; -- -0.025637604296207428
	pesos_i(2819) := b"0000000000000000_0000000000000000_0011001010000100_0001111110000000"; -- 0.19732853770256042
	pesos_i(2820) := b"0000000000000000_0000000000000000_0010111100001100_1100110011000000"; -- 0.18378905951976776
	pesos_i(2821) := b"0000000000000000_0000000000000000_0011111011110010_0000110010000000"; -- 0.2458808720111847
	pesos_i(2822) := b"0000000000000000_0000000000000000_0000010011011100_1011010111001000"; -- 0.018992768600583076
	pesos_i(2823) := b"1111111111111111_1111111111111111_1101100010011010_0000000101000000"; -- -0.15390007197856903
	pesos_i(2824) := b"1111111111111111_1111111111111111_1111101100111101_1010001011101000"; -- -0.01859075389802456
	pesos_i(2825) := b"0000000000000000_0000000000000000_0011011101010001_1010100000000000"; -- 0.21608972549438477
	pesos_i(2826) := b"0000000000000000_0000000000000000_0010000110010101_1010101101000000"; -- 0.13119001686573029
	pesos_i(2827) := b"1111111111111111_1111111111111111_1100011010001101_1110100001000000"; -- -0.22439716756343842
	pesos_i(2828) := b"1111111111111111_1111111111111111_1110101011010110_1010100111100000"; -- -0.08266199380159378
	pesos_i(2829) := b"1111111111111111_1111111111111111_1111111000000010_1101000111101000"; -- -0.007769471034407616
	pesos_i(2830) := b"1111111111111111_1111111111111111_1111100011110010_1110110110000000"; -- -0.027543216943740845
	pesos_i(2831) := b"0000000000000000_0000000000000000_0010000011001011_0001011000000000"; -- 0.12809884548187256
	pesos_i(2832) := b"1111111111111111_1111111111111111_1111010001011111_0110100011110000"; -- -0.04541916027665138
	pesos_i(2833) := b"0000000000000000_0000000000000000_0001101000010111_1000110100000000"; -- 0.10192185640335083
	pesos_i(2834) := b"1111111111111111_1111111111111111_1111100011100010_1100010000010000"; -- -0.027789827436208725
	pesos_i(2835) := b"1111111111111111_1111111111111111_1110110011111000_1101100010000000"; -- -0.07432791590690613
	pesos_i(2836) := b"0000000000000000_0000000000000000_0011010101001110_0011111000000000"; -- 0.20822513103485107
	pesos_i(2837) := b"1111111111111111_1111111111111111_1110000010011110_1111101000000000"; -- -0.12257421016693115
	pesos_i(2838) := b"0000000000000000_0000000000000000_0001101010100100_0111011011000000"; -- 0.10407201945781708
	pesos_i(2839) := b"1111111111111111_1111111111111111_1110101100110110_1011010010000000"; -- -0.08119651675224304
	pesos_i(2840) := b"0000000000000000_0000000000000000_0101000000010111_0000100100000000"; -- 0.3128514885902405
	pesos_i(2841) := b"1111111111111111_1111111111111111_1111111100110101_0010011101010100"; -- -0.003095190040767193
	pesos_i(2842) := b"1111111111111111_1111111111111111_1111011000110110_0001100000010000"; -- -0.03823709115386009
	pesos_i(2843) := b"0000000000000000_0000000000000000_0001010110110010_0001000011100000"; -- 0.08474832028150558
	pesos_i(2844) := b"0000000000000000_0000000000000000_0010011110101010_0001111100000000"; -- 0.15493959188461304
	pesos_i(2845) := b"0000000000000000_0000000000000000_0011101010110100_1101100001000000"; -- 0.22932197153568268
	pesos_i(2846) := b"0000000000000000_0000000000000000_0010100000101111_0011001101000000"; -- 0.15697021782398224
	pesos_i(2847) := b"1111111111111111_1111111111111111_1111111011010111_1000011101010110"; -- -0.004523793701082468
	pesos_i(2848) := b"0000000000000000_0000000000000000_0001001000010000_0101010100000000"; -- 0.07056170701980591
	pesos_i(2849) := b"1111111111111111_1111111111111111_1110110101111110_1100000010100000"; -- -0.07228466123342514
	pesos_i(2850) := b"0000000000000000_0000000000000000_0011111110011110_0000111000000000"; -- 0.24850547313690186
	pesos_i(2851) := b"0000000000000000_0000000000000000_0010101110110111_1100101000000000"; -- 0.17077314853668213
	pesos_i(2852) := b"1111111111111111_1111111111111111_1110111111101101_0011001100000000"; -- -0.06278687715530396
	pesos_i(2853) := b"0000000000000000_0000000000000000_0010100000011001_0010000010000000"; -- 0.1566334068775177
	pesos_i(2854) := b"0000000000000000_0000000000000000_0000000110011001_0010010110001100"; -- 0.006243082694709301
	pesos_i(2855) := b"1111111111111111_1111111111111111_1111101111110100_1010100111110000"; -- -0.015797976404428482
	pesos_i(2856) := b"0000000000000000_0000000000000000_0010000100100111_1111111010000000"; -- 0.12951651215553284
	pesos_i(2857) := b"1111111111111111_1111111111111111_1110110010001101_1101100101000000"; -- -0.07596056163311005
	pesos_i(2858) := b"0000000000000000_0000000000000000_0000010100000001_0001000100101000"; -- 0.019547531381249428
	pesos_i(2859) := b"1111111111111111_1111111111111111_1100101001100000_1100110100000000"; -- -0.20946043729782104
	pesos_i(2860) := b"1111111111111111_1111111111111111_1011011010000101_0011001010000000"; -- -0.28703007102012634
	pesos_i(2861) := b"0000000000000000_0000000000000000_0001110001100100_0001011010100000"; -- 0.11090222746133804
	pesos_i(2862) := b"0000000000000000_0000000000000000_0011001000111101_1111000110000000"; -- 0.19625768065452576
	pesos_i(2863) := b"0000000000000000_0000000000000000_0000101111000010_0000100111110000"; -- 0.045929547399282455
	pesos_i(2864) := b"0000000000000000_0000000000000000_0001100011010011_0000001111100000"; -- 0.096969835460186
	pesos_i(2865) := b"1111111111111111_1111111111111111_1010100011011101_0000100100000000"; -- -0.3403772711753845
	pesos_i(2866) := b"0000000000000000_0000000000000000_0000110101010110_0100011010010000"; -- 0.052097711712121964
	pesos_i(2867) := b"1111111111111111_1111111111111110_1110111101100111_1010111000000000"; -- -1.0648242235183716
	pesos_i(2868) := b"0000000000000000_0000000000000000_0001101011000000_0110001000100000"; -- 0.10449803620576859
	pesos_i(2869) := b"0000000000000000_0000000000000000_0001110010111101_0011010001100000"; -- 0.11226203292608261
	pesos_i(2870) := b"0000000000000000_0000000000000000_0011011000001101_0111111010000000"; -- 0.2111434042453766
	pesos_i(2871) := b"0000000000000000_0000000000000000_0000111010010001_0111001101000000"; -- 0.056906893849372864
	pesos_i(2872) := b"0000000000000000_0000000000000000_0010011001100110_0100100100000000"; -- 0.1499982476234436
	pesos_i(2873) := b"1111111111111111_1111111111111111_1100111101001111_1111101111000000"; -- -0.1901858001947403
	pesos_i(2874) := b"0000000000000000_0000000000000000_0000111111000110_1111001010000000"; -- 0.06162944436073303
	pesos_i(2875) := b"1111111111111111_1111111111111111_1111110011010110_1001011000100100"; -- -0.01235067006200552
	pesos_i(2876) := b"1111111111111111_1111111111111111_1111000010100111_0111010000100000"; -- -0.05994486063718796
	pesos_i(2877) := b"0000000000000000_0000000000000000_0001101011101100_0011001000100000"; -- 0.10516656190156937
	pesos_i(2878) := b"0000000000000000_0000000000000000_0001011011101001_1101111011100000"; -- 0.08950608223676682
	pesos_i(2879) := b"1111111111111111_1111111111111111_1000101111000100_0100111100000000"; -- -0.45403581857681274
	pesos_i(2880) := b"0000000000000000_0000000000000000_0100101101010110_1100101110000000"; -- 0.2942931354045868
	pesos_i(2881) := b"0000000000000000_0000000000000000_0010111101000111_1110101100000000"; -- 0.18469113111495972
	pesos_i(2882) := b"0000000000000000_0000000000000000_0000111100100000_0110101000010000"; -- 0.05908835306763649
	pesos_i(2883) := b"0000000000000000_0000000000000000_0011000011111110_1101100100000000"; -- 0.19138866662979126
	pesos_i(2884) := b"1111111111111111_1111111111111111_1110010011100100_1111010000100000"; -- -0.10588144510984421
	pesos_i(2885) := b"0000000000000000_0000000000000000_0000000010000000_1110010111101110"; -- 0.001966829877346754
	pesos_i(2886) := b"0000000000000000_0000000000000000_0101010000100111_1010100000000000"; -- 0.32873010635375977
	pesos_i(2887) := b"0000000000000000_0000000000000000_0000111000110001_1010100100110000"; -- 0.055445265024900436
	pesos_i(2888) := b"1111111111111111_1111111111111111_1111101101110001_0000000000100000"; -- -0.017806999385356903
	pesos_i(2889) := b"0000000000000000_0000000000000000_0000001011101001_0111100100110000"; -- 0.011375021189451218
	pesos_i(2890) := b"1111111111111111_1111111111111111_1011100111001101_1111010100000000"; -- -0.27420109510421753
	pesos_i(2891) := b"1111111111111111_1111111111111111_1101111100010000_0011001101000000"; -- -0.12865905463695526
	pesos_i(2892) := b"0000000000000000_0000000000000000_0001111010000111_0010110011000000"; -- 0.1192501038312912
	pesos_i(2893) := b"0000000000000000_0000000000000000_0010010101111011_1001110001000000"; -- 0.14641739428043365
	pesos_i(2894) := b"0000000000000000_0000000000000000_0001010010011110_0100110001100000"; -- 0.08054044097661972
	pesos_i(2895) := b"1111111111111111_1111111111111111_1101010000111110_1001100100000000"; -- -0.17091983556747437
	pesos_i(2896) := b"1111111111111111_1111111111111111_1101011001110011_1101000110000000"; -- -0.16229525208473206
	pesos_i(2897) := b"1111111111111111_1111111111111111_1011000000010111_0101010000000000"; -- -0.31214404106140137
	pesos_i(2898) := b"1111111111111111_1111111111111111_1110101000111110_1001011010000000"; -- -0.0849824845790863
	pesos_i(2899) := b"0000000000000000_0000000000000000_0001000100111001_1010101111100000"; -- 0.06728624552488327
	pesos_i(2900) := b"0000000000000000_0000000000000000_0001111110010010_1101100100100000"; -- 0.12333447486162186
	pesos_i(2901) := b"0000000000000000_0000000000000000_0100011111110000_0110110110000000"; -- 0.2810123860836029
	pesos_i(2902) := b"1111111111111111_1111111111111111_1111001101111011_0011010110010000"; -- -0.04890122637152672
	pesos_i(2903) := b"0000000000000000_0000000000000000_0011010111110100_0101101111000000"; -- 0.21075986325740814
	pesos_i(2904) := b"1111111111111111_1111111111111111_1100010101111100_0110000000000000"; -- -0.22857093811035156
	pesos_i(2905) := b"1111111111111111_1111111111111111_1110010110011011_0101100111100000"; -- -0.10309828072786331
	pesos_i(2906) := b"1111111111111111_1111111111111111_1101010110100010_0111100010000000"; -- -0.16548964381217957
	pesos_i(2907) := b"1111111111111111_1111111111111111_1111100111100110_0001101011110000"; -- -0.023832622915506363
	pesos_i(2908) := b"0000000000000000_0000000000000000_0001001001110010_1010100000000000"; -- 0.07206201553344727
	pesos_i(2909) := b"0000000000000000_0000000000000000_0011001011100001_0000100011000000"; -- 0.19874624907970428
	pesos_i(2910) := b"0000000000000000_0000000000000000_0000110111010101_0000010101110000"; -- 0.054031696170568466
	pesos_i(2911) := b"1111111111111111_1111111111111111_1110101110010001_1111100000100000"; -- -0.0798039361834526
	pesos_i(2912) := b"0000000000000000_0000000000000000_0011001011101000_0110011100000000"; -- 0.19885867834091187
	pesos_i(2913) := b"1111111111111111_1111111111111111_1110101010001100_0010100101000000"; -- -0.08379881083965302
	pesos_i(2914) := b"0000000000000000_0000000000000000_0010111100001101_0111010101000000"; -- 0.18379910290241241
	pesos_i(2915) := b"1111111111111111_1111111111111111_1111100111001000_0101110100101000"; -- -0.024286439642310143
	pesos_i(2916) := b"0000000000000000_0000000000000000_0000101100111010_0100011000010000"; -- 0.043857935816049576
	pesos_i(2917) := b"0000000000000000_0000000000000000_0010100011001110_0010001110000000"; -- 0.15939542651176453
	pesos_i(2918) := b"0000000000000000_0000000000000000_0000010001000111_0001011111011000"; -- 0.016709795221686363
	pesos_i(2919) := b"0000000000000000_0000000000000000_0011010100101110_1010111010000000"; -- 0.2077435553073883
	pesos_i(2920) := b"1111111111111111_1111111111111111_1111010101000000_1000010001010000"; -- -0.041984301060438156
	pesos_i(2921) := b"0000000000000000_0000000000000000_0001110001000011_1110111110000000"; -- 0.1104116141796112
	pesos_i(2922) := b"0000000000000000_0000000000000000_0000011101111111_1101001001111000"; -- 0.02929416112601757
	pesos_i(2923) := b"1111111111111111_1111111111111111_1111111111001000_0100100001111010"; -- -0.0008501723641529679
	pesos_i(2924) := b"1111111111111111_1111111111111111_0111100010010001_0001100100000000"; -- -0.5290359854698181
	pesos_i(2925) := b"0000000000000000_0000000000000000_0010000010101000_1111111000000000"; -- 0.12757861614227295
	pesos_i(2926) := b"1111111111111111_1111111111111111_1111000001010000_1001001100000000"; -- -0.06127053499221802
	pesos_i(2927) := b"1111111111111111_1111111111111111_1101111010001011_1000100001000000"; -- -0.13068340718746185
	pesos_i(2928) := b"1111111111111111_1111111111111111_1101100110111001_0011100101000000"; -- -0.1495174616575241
	pesos_i(2929) := b"0000000000000000_0000000000000000_0001111011101001_1011110100000000"; -- 0.12075406312942505
	pesos_i(2930) := b"1111111111111111_1111111111111111_1100110000010110_0110101000000000"; -- -0.2027829885482788
	pesos_i(2931) := b"1111111111111111_1111111111111111_1111000100111100_0100000001000000"; -- -0.05767439305782318
	pesos_i(2932) := b"0000000000000000_0000000000000000_0000101110101100_1100011111000000"; -- 0.045605167746543884
	pesos_i(2933) := b"1111111111111111_1111111111111111_1110111101110001_1011011000000000"; -- -0.06467115879058838
	pesos_i(2934) := b"0000000000000000_0000000000000000_0000101101110101_1101011011000000"; -- 0.044766828417778015
	pesos_i(2935) := b"0000000000000000_0000000000000000_0010001110111110_1001111000000000"; -- 0.1396273374557495
	pesos_i(2936) := b"1111111111111111_1111111111111111_1110001110101000_1011101100100000"; -- -0.1107066199183464
	pesos_i(2937) := b"0000000000000000_0000000000000000_0000000001110011_0001101101011000"; -- 0.001756390556693077
	pesos_i(2938) := b"1111111111111111_1111111111111111_1100101101011001_1100011101000000"; -- -0.205661341547966
	pesos_i(2939) := b"1111111111111111_1111111111111111_1110101011000101_0010111011000000"; -- -0.08292873203754425
	pesos_i(2940) := b"1111111111111111_1111111111111111_1111001010011101_0101101101000000"; -- -0.052286431193351746
	pesos_i(2941) := b"1111111111111111_1111111111111111_1101111101111000_0000000010000000"; -- -0.1270751655101776
	pesos_i(2942) := b"0000000000000000_0000000000000000_0001001111100101_1100001100000000"; -- 0.0777246356010437
	pesos_i(2943) := b"0000000000000000_0000000000000000_0000111001011111_0110010001100000"; -- 0.05614306777715683
	pesos_i(2944) := b"1111111111111111_1111111111111111_1110101111010110_1001010001100000"; -- -0.07875702530145645
	pesos_i(2945) := b"0000000000000000_0000000000000000_0000011110000001_1111011100011000"; -- 0.02932686172425747
	pesos_i(2946) := b"1111111111111111_1111111111111111_1101011101010110_0111111110000000"; -- -0.15883639454841614
	pesos_i(2947) := b"0000000000000000_0000000000000000_0111110100101011_0010110110000000"; -- 0.4889400899410248
	pesos_i(2948) := b"1111111111111111_1111111111111111_1101011010111110_1100110100000000"; -- -0.16115111112594604
	pesos_i(2949) := b"0000000000000000_0000000000000000_0011100010010010_0101111111000000"; -- 0.22098349034786224
	pesos_i(2950) := b"1111111111111111_1111111111111111_1110101101111101_1011001011000000"; -- -0.0801132470369339
	pesos_i(2951) := b"0000000000000000_0000000000000000_0001001010110100_0011110011000000"; -- 0.0730627030134201
	pesos_i(2952) := b"1111111111111111_1111111111111111_1110000100110101_1000000001000000"; -- -0.12027738988399506
	pesos_i(2953) := b"0000000000000000_0000000000000000_0101010001000011_1111011010000000"; -- 0.32916203141212463
	pesos_i(2954) := b"1111111111111111_1111111111111111_1110000011011110_0111010111100000"; -- -0.1216055229306221
	pesos_i(2955) := b"1111111111111111_1111111111111111_1101011111001011_1010001011000000"; -- -0.1570490151643753
	pesos_i(2956) := b"0000000000000000_0000000000000000_0011000000001011_0000101110000000"; -- 0.18766853213310242
	pesos_i(2957) := b"0000000000000000_0000000000000000_0001011110010101_1101111110100000"; -- 0.0921306386590004
	pesos_i(2958) := b"1111111111111111_1111111111111111_1100110101101101_1011111100000000"; -- -0.1975441575050354
	pesos_i(2959) := b"1111111111111111_1111111111111111_1110000000111000_1100010110000000"; -- -0.12413373589515686
	pesos_i(2960) := b"1111111111111111_1111111111111111_1111001011100111_1100010111110000"; -- -0.05115092173218727
	pesos_i(2961) := b"1111111111111111_1111111111111111_1110110101111110_1011101101100000"; -- -0.07228497415781021
	pesos_i(2962) := b"0000000000000000_0000000000000000_0001001000110100_0011001100100000"; -- 0.07110900431871414
	pesos_i(2963) := b"1111111111111111_1111111111111111_1101101111100010_1101001011000000"; -- -0.1410702019929886
	pesos_i(2964) := b"0000000000000000_0000000000000000_0010110011001111_1110100100000000"; -- 0.17504745721817017
	pesos_i(2965) := b"1111111111111111_1111111111111111_1101110000111001_0001111111000000"; -- -0.13975335657596588
	pesos_i(2966) := b"1111111111111111_1111111111111111_1111001101100000_1010011001110000"; -- -0.049306485801935196
	pesos_i(2967) := b"1111111111111111_1111111111111111_1101101011100000_0001010100000000"; -- -0.14501827955245972
	pesos_i(2968) := b"0000000000000000_0000000000000000_0010001011010100_0110011100000000"; -- 0.13605350255966187
	pesos_i(2969) := b"0000000000000000_0000000000000000_0100110100011010_0001001010000000"; -- 0.30117908120155334
	pesos_i(2970) := b"1111111111111111_1111111111111111_1000011001011000_1101000110000000"; -- -0.47520723938941956
	pesos_i(2971) := b"1111111111111111_1111111111111111_1111101000000101_1100101001001000"; -- -0.023349149152636528
	pesos_i(2972) := b"0000000000000000_0000000000000000_0001111101110011_1010000001000000"; -- 0.12285806238651276
	pesos_i(2973) := b"0000000000000000_0000000000000000_0011010100010011_0111011111000000"; -- 0.20732830464839935
	pesos_i(2974) := b"1111111111111111_1111111111111111_1100111000001111_1010101110000000"; -- -0.19507339596748352
	pesos_i(2975) := b"0000000000000000_0000000000000000_0001001100101010_1001110101100000"; -- 0.07486899942159653
	pesos_i(2976) := b"0000000000000000_0000000000000000_0001111011111011_0010011100100000"; -- 0.12101978808641434
	pesos_i(2977) := b"1111111111111111_1111111111111111_1101011001000101_1011111111000000"; -- -0.16299821436405182
	pesos_i(2978) := b"0000000000000000_0000000000000000_0101101001011000_0110100100000000"; -- 0.3529115319252014
	pesos_i(2979) := b"0000000000000000_0000000000000000_0100100101100100_0100000100000000"; -- 0.2866860032081604
	pesos_i(2980) := b"0000000000000000_0000000000000000_0011110010111110_0111101111000000"; -- 0.23728154599666595
	pesos_i(2981) := b"0000000000000000_0000000000000000_0000100011101111_0010010111110000"; -- 0.034899111837148666
	pesos_i(2982) := b"1111111111111111_1111111111111111_1101111100100000_0110001010000000"; -- -0.12841209769248962
	pesos_i(2983) := b"0000000000000000_0000000000000000_0001001101001011_1000011111100000"; -- 0.07537125796079636
	pesos_i(2984) := b"0000000000000000_0000000000000000_0001110100010010_1110101001100000"; -- 0.11356987804174423
	pesos_i(2985) := b"1111111111111111_1111111111111111_1110100000111110_1000010101100000"; -- -0.09279600530862808
	pesos_i(2986) := b"0000000000000000_0000000000000000_0001010001100010_1011110100100000"; -- 0.07963163405656815
	pesos_i(2987) := b"1111111111111111_1111111111111111_1010111001010101_0100010000000000"; -- -0.3190114498138428
	pesos_i(2988) := b"1111111111111111_1111111111111111_1101100000111101_0110110010000000"; -- -0.15531274676322937
	pesos_i(2989) := b"1111111111111111_1111111111111111_1110100000100001_1110000110100000"; -- -0.09323301166296005
	pesos_i(2990) := b"0000000000000000_0000000000000000_0000001000001011_0100011111001100"; -- 0.007984626106917858
	pesos_i(2991) := b"0000000000000000_0000000000000000_0010100011001000_1100000101000000"; -- 0.15931327641010284
	pesos_i(2992) := b"0000000000000000_0000000000000000_0011111000001101_1101100101000000"; -- 0.24239881336688995
	pesos_i(2993) := b"1111111111111111_1111111111111111_1101000100101100_1101010110000000"; -- -0.18290963768959045
	pesos_i(2994) := b"1111111111111111_1111111111111111_1101100010000101_1010011110000000"; -- -0.15421059727668762
	pesos_i(2995) := b"1111111111111111_1111111111111111_1001100101110110_1001100000000000"; -- -0.40053415298461914
	pesos_i(2996) := b"0000000000000000_0000000000000000_0010111111000101_1011001100000000"; -- 0.1866104006767273
	pesos_i(2997) := b"0000000000000000_0000000000000000_0010010100001011_1110100000000000"; -- 0.1447129249572754
	pesos_i(2998) := b"0000000000000000_0000000000000000_0011000010110000_1101000000000000"; -- 0.19019794464111328
	pesos_i(2999) := b"1111111111111111_1111111111111111_1111000111011000_1110101101000000"; -- -0.05528382956981659
	pesos_i(3000) := b"0000000000000000_0000000000000000_0100010011100111_1101110110000000"; -- 0.26916298270225525
	pesos_i(3001) := b"1111111111111111_1111111111111111_1101100000001010_1110110011000000"; -- -0.15608330070972443
	pesos_i(3002) := b"1111111111111111_1111111111111111_1110100011011011_0111000001100000"; -- -0.09040162712335587
	pesos_i(3003) := b"0000000000000000_0000000000000000_0000001110111011_0011101000011100"; -- 0.014575607143342495
	pesos_i(3004) := b"0000000000000000_0000000000000000_0001011110111111_1100011010000000"; -- 0.09277001023292542
	pesos_i(3005) := b"1111111111111111_1111111111111111_1111001100000100_0100001100100000"; -- -0.05071621388196945
	pesos_i(3006) := b"1111111111111111_1111111111111111_1111000001001011_0100000100100000"; -- -0.0613517090678215
	pesos_i(3007) := b"1111111111111111_1111111111111111_1000111101111101_0011111100000000"; -- -0.43949514627456665
	pesos_i(3008) := b"0000000000000000_0000000000000000_0000011110010001_0110110011111000"; -- 0.02956276945769787
	pesos_i(3009) := b"0000000000000000_0000000000000000_0010110010101001_0011000100000000"; -- 0.1744566559791565
	pesos_i(3010) := b"0000000000000000_0000000000000000_0010011010000011_0000101000000000"; -- 0.15043699741363525
	pesos_i(3011) := b"0000000000000000_0000000000000000_0000000110101000_1010011011111000"; -- 0.006479678675532341
	pesos_i(3012) := b"1111111111111111_1111111111111111_1001100111111001_0100000100000000"; -- -0.3985404372215271
	pesos_i(3013) := b"0000000000000000_0000000000000000_0000001110001001_0100010100101100"; -- 0.013813327066600323
	pesos_i(3014) := b"0000000000000000_0000000000000000_0011001100011010_1100000000000000"; -- 0.19962692260742188
	pesos_i(3015) := b"1111111111111111_1111111111111111_1111010111100000_1010111001000000"; -- -0.03954039514064789
	pesos_i(3016) := b"0000000000000000_0000000000000000_0001111011001011_0000100111100000"; -- 0.12028562277555466
	pesos_i(3017) := b"1111111111111111_1111111111111111_1111110000101000_1010000001000100"; -- -0.015005095861852169
	pesos_i(3018) := b"1111111111111111_1111111111111111_1100110000111001_0011011110000000"; -- -0.20225194096565247
	pesos_i(3019) := b"0000000000000000_0000000000000000_0000111010010111_1010100111110000"; -- 0.05700170621275902
	pesos_i(3020) := b"0000000000000000_0000000000000000_0001101000001101_1101101010000000"; -- 0.10177388787269592
	pesos_i(3021) := b"1111111111111111_1111111111111111_1101001111111101_1111110011000000"; -- -0.17190571129322052
	pesos_i(3022) := b"1111111111111111_1111111111111111_1110000011100011_0000110111000000"; -- -0.12153543531894684
	pesos_i(3023) := b"1111111111111111_1111111111111111_1011000110110101_1001001010000000"; -- -0.3058231770992279
	pesos_i(3024) := b"1111111111111111_1111111111111111_1110100010001101_1001101111100000"; -- -0.09158921986818314
	pesos_i(3025) := b"1111111111111111_1111111111111111_0111100001111011_1010000100000000"; -- -0.5293635725975037
	pesos_i(3026) := b"0000000000000000_0000000000000000_0010110111110101_0101111111000000"; -- 0.17952536046504974
	pesos_i(3027) := b"0000000000000000_0000000000000000_0010101001110101_0101111111000000"; -- 0.16585348546504974
	pesos_i(3028) := b"0000000000000000_0000000000000000_0110001101110101_0011001000000000"; -- 0.38850700855255127
	pesos_i(3029) := b"0000000000000000_0000000000000000_0010100110100001_0101100011000000"; -- 0.16261820495128632
	pesos_i(3030) := b"1111111111111111_1111111111111111_1111000011110000_0110011101000000"; -- -0.05883173644542694
	pesos_i(3031) := b"0000000000000000_0000000000000000_0001100001000011_0010001000000000"; -- 0.09477436542510986
	pesos_i(3032) := b"1111111111111111_1111111111111111_1010010101111010_1001001110000000"; -- -0.35359838604927063
	pesos_i(3033) := b"0000000000000000_0000000000000000_0101001011001100_0110010100000000"; -- 0.3234313130378723
	pesos_i(3034) := b"1111111111111111_1111111111111111_1100011111111010_0111110100000000"; -- -0.21883410215377808
	pesos_i(3035) := b"1111111111111111_1111111111111111_1010011101100101_0111100100000000"; -- -0.3461079001426697
	pesos_i(3036) := b"0000000000000000_0000000000000000_0000110010100101_1100101010110000"; -- 0.04940478131175041
	pesos_i(3037) := b"0000000000000000_0000000000000000_0000001101111110_1001001111010000"; -- 0.013650167733430862
	pesos_i(3038) := b"1111111111111111_1111111111111111_1111010011000110_0010001010010000"; -- -0.04385169968008995
	pesos_i(3039) := b"1111111111111111_1111111111111111_1001001011001000_1000100010000000"; -- -0.42662760615348816
	pesos_i(3040) := b"0000000000000000_0000000000000000_0010011001001001_0110110110000000"; -- 0.1495579183101654
	pesos_i(3041) := b"0000000000000000_0000000000000000_0000010011100011_1000010110001000"; -- 0.019096704199910164
	pesos_i(3042) := b"1111111111111111_1111111111111111_1111001010110110_1111100100000000"; -- -0.05189555883407593
	pesos_i(3043) := b"1111111111111111_1111111111111111_1100100000101110_0110000110000000"; -- -0.2180422842502594
	pesos_i(3044) := b"1111111111111111_1111111111111111_1111010101010111_0010011110010000"; -- -0.041638877242803574
	pesos_i(3045) := b"0000000000000000_0000000000000000_0000101011000110_0101111110010000"; -- 0.04208943620324135
	pesos_i(3046) := b"0000000000000000_0000000000000000_0001101111010001_0001111111000000"; -- 0.10865972936153412
	pesos_i(3047) := b"1111111111111111_1111111111111111_1110101100110011_0011101000000000"; -- -0.08124959468841553
	pesos_i(3048) := b"0000000000000000_0000000000000000_0001000011101100_1110100001000000"; -- 0.06611491739749908
	pesos_i(3049) := b"0000000000000000_0000000000000000_0001100111110000_1001010000000000"; -- 0.10132718086242676
	pesos_i(3050) := b"1111111111111111_1111111111111111_1111001100101011_0101111101010000"; -- -0.050119441002607346
	pesos_i(3051) := b"0000000000000000_0000000000000000_0000111011011011_1001110110110000"; -- 0.05803857371211052
	pesos_i(3052) := b"1111111111111111_1111111111111111_1100010011001101_0011001100000000"; -- -0.23124390840530396
	pesos_i(3053) := b"0000000000000000_0000000000000000_0000001001111111_1100101010100100"; -- 0.009762444533407688
	pesos_i(3054) := b"1111111111111111_1111111111111111_1110000111000101_1011011101000000"; -- -0.11807684600353241
	pesos_i(3055) := b"0000000000000000_0000000000000000_0000101000000101_0111010000110000"; -- 0.03914571925997734
	pesos_i(3056) := b"0000000000000000_0000000000000000_0010011110101010_1111000100000000"; -- 0.15495210886001587
	pesos_i(3057) := b"0000000000000000_0000000000000000_0011000100011101_1001010111000000"; -- 0.19185768067836761
	pesos_i(3058) := b"1111111111111111_1111111111111111_1110001001000000_0111101101100000"; -- -0.11620358377695084
	pesos_i(3059) := b"1111111111111111_1111111111111111_1110011000011000_0111011000000000"; -- -0.1011892557144165
	pesos_i(3060) := b"0000000000000000_0000000000000000_0100000110111100_1001100000000000"; -- 0.25678396224975586
	pesos_i(3061) := b"1111111111111111_1111111111111111_1001110011011110_0111010100000000"; -- -0.3872305750846863
	pesos_i(3062) := b"1111111111111111_1111111111111111_1010001111000111_0000000110000000"; -- -0.36024466156959534
	pesos_i(3063) := b"1111111111111111_1111111111111111_1001111110101000_1011011010000000"; -- -0.3763318955898285
	pesos_i(3064) := b"1111111111111111_1111111111111111_1111100000101001_1000000111010000"; -- -0.030616652220487595
	pesos_i(3065) := b"1111111111111111_1111111111111111_1110001000000100_0110111111000000"; -- -0.11711980402469635
	pesos_i(3066) := b"1111111111111111_1111111111111111_1111100110100101_1101100011010000"; -- -0.024813126772642136
	pesos_i(3067) := b"0000000000000000_0000000000000000_0001000001101111_1010011100000000"; -- 0.06420367956161499
	pesos_i(3068) := b"0000000000000000_0000000000000000_0000110110110101_0111100100010000"; -- 0.05355030670762062
	pesos_i(3069) := b"1111111111111111_1111111111111111_1100001000000010_1100101101000000"; -- -0.2421448677778244
	pesos_i(3070) := b"0000000000000000_0000000000000000_0100001111011111_1000110100000000"; -- 0.26512986421585083
	pesos_i(3071) := b"1111111111111111_1111111111111111_1100000001010100_0100111100000000"; -- -0.24871355295181274
	pesos_i(3072) := b"0000000000000000_0000000000000000_0001010110100000_0000101110000000"; -- 0.08447334170341492
	pesos_i(3073) := b"0000000000000000_0000000000000000_0011101011100111_0100110100000000"; -- 0.2300918698310852
	pesos_i(3074) := b"1111111111111111_1111111111111111_1111011010001100_1110010100000000"; -- -0.036912620067596436
	pesos_i(3075) := b"1111111111111111_1111111111111111_1101100110101001_1011010100000000"; -- -0.14975422620773315
	pesos_i(3076) := b"0000000000000000_0000000000000000_0010001011100101_1111101101000000"; -- 0.13632173836231232
	pesos_i(3077) := b"1111111111111111_1111111111111111_1101001101111100_0110110101000000"; -- -0.1738826483488083
	pesos_i(3078) := b"1111111111111111_1111111111111111_1110100001100100_0100001011100000"; -- -0.09222013503313065
	pesos_i(3079) := b"0000000000000000_0000000000000000_0000111011011000_1000101010010000"; -- 0.05799165740609169
	pesos_i(3080) := b"0000000000000000_0000000000000000_0001000010000100_1110100001000000"; -- 0.06452800333499908
	pesos_i(3081) := b"1111111111111111_1111111111111111_1100011101000101_0110011100000000"; -- -0.22159725427627563
	pesos_i(3082) := b"0000000000000000_0000000000000000_0011100111000010_1000000100000000"; -- 0.22562414407730103
	pesos_i(3083) := b"0000000000000000_0000000000000000_0100010011010110_0110001110000000"; -- 0.26889631152153015
	pesos_i(3084) := b"1111111111111111_1111111111111111_1111100111111100_1100101010100000"; -- -0.023486457765102386
	pesos_i(3085) := b"1111111111111111_1111111111111111_1010111001110011_1010100000000000"; -- -0.31854772567749023
	pesos_i(3086) := b"0000000000000000_0000000000000000_0001000110111000_1001000111000000"; -- 0.06922255456447601
	pesos_i(3087) := b"0000000000000000_0000000000000000_0000010101001001_1101101100101000"; -- 0.020658204331994057
	pesos_i(3088) := b"1111111111111111_1111111111111111_1100011010100100_1000000101000000"; -- -0.22405235469341278
	pesos_i(3089) := b"0000000000000000_0000000000000000_0000010011101110_0001100101111000"; -- 0.019258109852671623
	pesos_i(3090) := b"0000000000000000_0000000000000000_0010011110000010_1000100100000000"; -- 0.15433555841445923
	pesos_i(3091) := b"0000000000000000_0000000000000000_0000110010010111_1100110100010000"; -- 0.049191299825906754
	pesos_i(3092) := b"1111111111111111_1111111111111111_1111111111010100_1101001011101100"; -- -0.0006588147953152657
	pesos_i(3093) := b"1111111111111111_1111111111111111_1110000001101101_0110100111100000"; -- -0.1233304813504219
	pesos_i(3094) := b"0000000000000000_0000000000000000_0001111010110110_1011011011100000"; -- 0.1199754998087883
	pesos_i(3095) := b"1111111111111111_1111111111111111_1101000110001011_0101101100000000"; -- -0.18146735429763794
	pesos_i(3096) := b"1111111111111111_1111111111111111_1100101101011110_1111000110000000"; -- -0.20558252930641174
	pesos_i(3097) := b"0000000000000000_0000000000000000_0000010110000011_0100000110100000"; -- 0.021534062922000885
	pesos_i(3098) := b"0000000000000000_0000000000000000_0010001010101000_1011001101000000"; -- 0.135386660695076
	pesos_i(3099) := b"1111111111111111_1111111111111111_1101100110001110_0000101101000000"; -- -0.15017633140087128
	pesos_i(3100) := b"0000000000000000_0000000000000000_0010111100011101_0010011001000000"; -- 0.18403853476047516
	pesos_i(3101) := b"1111111111111111_1111111111111111_1100011011111110_1101100100000000"; -- -0.22267383337020874
	pesos_i(3102) := b"0000000000000000_0000000000000000_0010000011110001_0110010001000000"; -- 0.12868334352970123
	pesos_i(3103) := b"1111111111111111_1111111111111111_1111011111011011_0000001101010000"; -- -0.03181437775492668
	pesos_i(3104) := b"0000000000000000_0000000000000000_0000111011001110_1011111101100000"; -- 0.05784221738576889
	pesos_i(3105) := b"0000000000000000_0000000000000000_0100011100110100_1010010010000000"; -- 0.27814701199531555
	pesos_i(3106) := b"0000000000000000_0000000000000000_0000101100110101_1000001100100000"; -- 0.04378528147935867
	pesos_i(3107) := b"0000000000000000_0000000000000000_0000000100110011_1100111001110000"; -- 0.00469675287604332
	pesos_i(3108) := b"1111111111111111_1111111111111111_1110111110010100_1110101011000000"; -- -0.06413395702838898
	pesos_i(3109) := b"1111111111111111_1111111111111111_1110010001100110_1001111110100000"; -- -0.10780908912420273
	pesos_i(3110) := b"1111111111111111_1111111111111111_1011110001011110_0111100100000000"; -- -0.2641834616661072
	pesos_i(3111) := b"0000000000000000_0000000000000000_0010110101100101_1101111111000000"; -- 0.177335724234581
	pesos_i(3112) := b"0000000000000000_0000000000000000_0000010011111101_0011011100110000"; -- 0.019488763064146042
	pesos_i(3113) := b"1111111111111111_1111111111111111_1111001000101110_1110010000110000"; -- -0.053971994668245316
	pesos_i(3114) := b"0000000000000000_0000000000000000_0000100000001010_1001110011100000"; -- 0.03141193836927414
	pesos_i(3115) := b"0000000000000000_0000000000000000_0000000011100110_0111100111010110"; -- 0.003516783472150564
	pesos_i(3116) := b"1111111111111111_1111111111111111_1111010100010000_0101101000000000"; -- -0.042719244956970215
	pesos_i(3117) := b"1111111111111111_1111111111111111_1110010000100000_1011101011000000"; -- -0.1088755875825882
	pesos_i(3118) := b"1111111111111111_1111111111111111_1111101011111010_1011101100100000"; -- -0.019611649215221405
	pesos_i(3119) := b"1111111111111111_1111111111111111_1110001101000010_0010101111000000"; -- -0.11227156221866608
	pesos_i(3120) := b"1111111111111111_1111111111111111_1110001111110101_0101110011000000"; -- -0.10953731834888458
	pesos_i(3121) := b"1111111111111111_1111111111111111_1101001001001010_0101001110000000"; -- -0.17855337262153625
	pesos_i(3122) := b"1111111111111111_1111111111111111_1000100010000011_0011011110000000"; -- -0.46674779057502747
	pesos_i(3123) := b"0000000000000000_0000000000000000_0011101111101110_1000111001000000"; -- 0.2341088205575943
	pesos_i(3124) := b"1111111111111111_1111111111111111_1110100010000010_0000011010100000"; -- -0.09176596254110336
	pesos_i(3125) := b"1111111111111111_1111111111111111_1111110111110010_0000010101111000"; -- -0.008025797083973885
	pesos_i(3126) := b"0000000000000000_0000000000000000_0000011110100011_0000000011011000"; -- 0.02983098290860653
	pesos_i(3127) := b"1111111111111111_1111111111111111_1111010000111010_0000011001100000"; -- -0.04598961025476456
	pesos_i(3128) := b"1111111111111111_1111111111111111_1100000110100100_0010100101000000"; -- -0.24358884990215302
	pesos_i(3129) := b"0000000000000000_0000000000000000_0010100101011101_0100011000000000"; -- 0.16157948970794678
	pesos_i(3130) := b"0000000000000000_0000000000000000_0010000111000011_1101111110000000"; -- 0.1318950355052948
	pesos_i(3131) := b"0000000000000000_0000000000000000_0000100101101011_1100110111010000"; -- 0.036801207810640335
	pesos_i(3132) := b"0000000000000000_0000000000000000_0100101001100001_1001011000000000"; -- 0.2905515432357788
	pesos_i(3133) := b"1111111111111111_1111111111111111_1111111011010101_0110100110011110"; -- -0.004556082654744387
	pesos_i(3134) := b"0000000000000000_0000000000000000_0001100001111111_0010101010100000"; -- 0.09569040685892105
	pesos_i(3135) := b"1111111111111111_1111111111111111_1100101101100110_0000100001000000"; -- -0.2054743617773056
	pesos_i(3136) := b"1111111111111111_1111111111111111_1101111010101111_0100000011000000"; -- -0.1301383525133133
	pesos_i(3137) := b"0000000000000000_0000000000000000_0011000000101111_0010010010000000"; -- 0.1882193386554718
	pesos_i(3138) := b"1111111111111111_1111111111111111_1101001101011000_1111110111000000"; -- -0.17442335188388824
	pesos_i(3139) := b"0000000000000000_0000000000000000_0010110100001110_1001011011000000"; -- 0.1760038584470749
	pesos_i(3140) := b"0000000000000000_0000000000000000_0001100100011001_1101010100000000"; -- 0.09805041551589966
	pesos_i(3141) := b"1111111111111111_1111111111111111_1111010111101101_1010110011010000"; -- -0.03934211656451225
	pesos_i(3142) := b"0000000000000000_0000000000000000_0011110111011010_0111101111000000"; -- 0.24161504209041595
	pesos_i(3143) := b"0000000000000000_0000000000000000_0001011101110001_1011111101000000"; -- 0.0915793925523758
	pesos_i(3144) := b"0000000000000000_0000000000000000_0010111111010111_1011000011000000"; -- 0.18688492476940155
	pesos_i(3145) := b"0000000000000000_0000000000000000_0010000011110010_1010010110000000"; -- 0.12870249152183533
	pesos_i(3146) := b"1111111111111111_1111111111111111_1111110001111000_0101001001000100"; -- -0.01378904189914465
	pesos_i(3147) := b"0000000000000000_0000000000000000_0011000001001000_0111100110000000"; -- 0.1886058747768402
	pesos_i(3148) := b"1111111111111111_1111111111111111_1110011110101011_0111100001000000"; -- -0.09503982961177826
	pesos_i(3149) := b"0000000000000000_0000000000000000_0100011101101101_1000010100000000"; -- 0.2790148854255676
	pesos_i(3150) := b"1111111111111111_1111111111111111_1010110111001011_0001001110000000"; -- -0.3211200535297394
	pesos_i(3151) := b"1111111111111111_1111111111111111_1111111010101101_1001100101010100"; -- -0.005163590423762798
	pesos_i(3152) := b"1111111111111111_1111111111111111_1100101111110100_1101100100000000"; -- -0.20329517126083374
	pesos_i(3153) := b"0000000000000000_0000000000000000_0001010010011111_0011001000100000"; -- 0.08055413514375687
	pesos_i(3154) := b"1111111111111111_1111111111111111_1011101000100011_0010100110000000"; -- -0.2729009687900543
	pesos_i(3155) := b"1111111111111111_1111111111111111_1110001111100111_1001001101000000"; -- -0.10974769294261932
	pesos_i(3156) := b"0000000000000000_0000000000000000_0010101011101011_0000100001000000"; -- 0.1676488071680069
	pesos_i(3157) := b"0000000000000000_0000000000000000_0011001111000101_1101010101000000"; -- 0.20223744213581085
	pesos_i(3158) := b"1111111111111111_1111111111111111_1101111010100011_0010110100000000"; -- -0.1303226351737976
	pesos_i(3159) := b"0000000000000000_0000000000000000_0000001110111101_0010100100111000"; -- 0.014605117961764336
	pesos_i(3160) := b"0000000000000000_0000000000000000_0000111110011101_1111011101000000"; -- 0.061004117131233215
	pesos_i(3161) := b"0000000000000000_0000000000000000_0001001100011011_1111000111100000"; -- 0.07464515417814255
	pesos_i(3162) := b"0000000000000000_0000000000000000_0000100010110100_1111100000100000"; -- 0.034011371433734894
	pesos_i(3163) := b"1111111111111111_1111111111111111_1100000001100101_1110010101000000"; -- -0.24844519793987274
	pesos_i(3164) := b"1111111111111111_1111111111111111_1010111011111000_0001001110000000"; -- -0.3165271580219269
	pesos_i(3165) := b"1111111111111111_1111111111111111_1101110110011101_0110101010000000"; -- -0.13431677222251892
	pesos_i(3166) := b"0000000000000000_0000000000000000_0010001110110100_0010010100000000"; -- 0.1394675374031067
	pesos_i(3167) := b"0000000000000000_0000000000000000_0011000111001110_1101101000000000"; -- 0.19456255435943604
	pesos_i(3168) := b"1111111111111111_1111111111111111_1110111111100000_1000011101000000"; -- -0.06298021972179413
	pesos_i(3169) := b"0000000000000000_0000000000000000_0000011110011110_1010111111000000"; -- 0.029765114188194275
	pesos_i(3170) := b"0000000000000000_0000000000000000_0110000111001000_1110100010000000"; -- 0.3819718658924103
	pesos_i(3171) := b"1111111111111111_1111111111111111_1101111010010011_0000100010000000"; -- -0.1305689513683319
	pesos_i(3172) := b"0000000000000000_0000000000000000_0010000100100011_1111101011000000"; -- 0.12945525348186493
	pesos_i(3173) := b"1111111111111111_1111111111111111_1111011010110011_1000010111010000"; -- -0.03632320091128349
	pesos_i(3174) := b"1111111111111111_1111111111111111_1110100100110010_0111100010000000"; -- -0.08907362818717957
	pesos_i(3175) := b"1111111111111111_1111111111111111_1010110001100111_0001000110000000"; -- -0.32655230164527893
	pesos_i(3176) := b"1111111111111111_1111111111111111_1101100111001100_0111001001000000"; -- -0.1492241472005844
	pesos_i(3177) := b"0000000000000000_0000000000000000_0010101010111001_1010111101000000"; -- 0.1668958216905594
	pesos_i(3178) := b"1111111111111111_1111111111111111_1110110100010100_1011111010100000"; -- -0.07390221208333969
	pesos_i(3179) := b"1111111111111111_1111111111111111_1111101000110111_0001100000000000"; -- -0.02259683609008789
	pesos_i(3180) := b"0000000000000000_0000000000000000_0001001000110111_0011110010100000"; -- 0.07115534693002701
	pesos_i(3181) := b"1111111111111111_1111111111111111_1000110000011110_0010110000000000"; -- -0.4526646137237549
	pesos_i(3182) := b"1111111111111111_1111111111111111_1111110001001001_0100000010000000"; -- -0.014507263898849487
	pesos_i(3183) := b"1111111111111111_1111111111111111_1101001100011110_1101111100000000"; -- -0.1753101944923401
	pesos_i(3184) := b"0000000000000000_0000000000000000_0000000111000110_1000000101001110"; -- 0.00693519739434123
	pesos_i(3185) := b"1111111111111111_1111111111111111_1010001000100101_1100000100000000"; -- -0.36661142110824585
	pesos_i(3186) := b"1111111111111111_1111111111111111_1111100010000001_1100010000010000"; -- -0.029269929975271225
	pesos_i(3187) := b"0000000000000000_0000000000000000_0011001001111110_0110110110000000"; -- 0.1972416341304779
	pesos_i(3188) := b"1111111111111111_1111111111111111_1110001110111001_0111000001000000"; -- -0.11045168340206146
	pesos_i(3189) := b"1111111111111111_1111111111111111_1101000000001010_1100000011000000"; -- -0.18733592331409454
	pesos_i(3190) := b"1111111111111111_1111111111111111_1111011011011110_1001001000000000"; -- -0.03566634654998779
	pesos_i(3191) := b"0000000000000000_0000000000000000_0010100010000010_1000011000000000"; -- 0.1582416296005249
	pesos_i(3192) := b"1111111111111111_1111111111111111_1101110100111010_0011100000000000"; -- -0.13583040237426758
	pesos_i(3193) := b"0000000000000000_0000000000000000_0001111100100010_0100011011000000"; -- 0.12161676585674286
	pesos_i(3194) := b"1111111111111111_1111111111111111_1101111110111111_0010011000000000"; -- -0.12598955631256104
	pesos_i(3195) := b"0000000000000000_0000000000000000_0010000001100011_1010100000000000"; -- 0.12652063369750977
	pesos_i(3196) := b"1111111111111111_1111111111111111_1101011100010101_0110101110000000"; -- -0.15982940793037415
	pesos_i(3197) := b"1111111111111111_1111111111111111_1101011100101111_0000001101000000"; -- -0.15943889319896698
	pesos_i(3198) := b"1111111111111111_1111111111111111_1101110010100111_0101110101000000"; -- -0.1380712240934372
	pesos_i(3199) := b"1111111111111111_1111111111111111_1110011110101101_1101110100100000"; -- -0.09500329941511154
	pesos_i(3200) := b"1111111111111111_1111111111111111_1101100001111100_1100001100000000"; -- -0.1543462872505188
	pesos_i(3201) := b"0000000000000000_0000000000000000_0100010011100001_0111010100000000"; -- 0.2690652012825012
	pesos_i(3202) := b"1111111111111111_1111111111111111_0111001100011101_0010100100000000"; -- -0.5503363013267517
	pesos_i(3203) := b"0000000000000000_0000000000000000_0001100011010101_0011100100100000"; -- 0.0970035269856453
	pesos_i(3204) := b"1111111111111111_1111111111111111_1111111001111001_0101111010100000"; -- -0.005960546433925629
	pesos_i(3205) := b"1111111111111111_1111111111111111_1011001010101111_0000111110000000"; -- -0.3020162880420685
	pesos_i(3206) := b"0000000000000000_0000000000000000_0010001001001011_1100010011000000"; -- 0.13396863639354706
	pesos_i(3207) := b"1111111111111111_1111111111111111_1111011011110101_1111010111000000"; -- -0.03530944883823395
	pesos_i(3208) := b"1111111111111111_1111111111111111_1111111011100001_1011111011101010"; -- -0.004367893096059561
	pesos_i(3209) := b"1111111111111111_1111111111111111_1110011011100110_1100101001100000"; -- -0.09804091602563858
	pesos_i(3210) := b"0000000000000000_0000000000000000_0010110100100100_0111001000000000"; -- 0.1763373613357544
	pesos_i(3211) := b"0000000000000000_0000000000000000_0001010010000110_0111111010000000"; -- 0.08017721772193909
	pesos_i(3212) := b"1111111111111111_1111111111111111_1111000001100011_0100110110000000"; -- -0.06098476052284241
	pesos_i(3213) := b"1111111111111111_1111111111111111_1100111011011111_0100101100000000"; -- -0.19190531969070435
	pesos_i(3214) := b"1111111111111111_1111111111111111_1001110101111100_0101011010000000"; -- -0.38482150435447693
	pesos_i(3215) := b"1111111111111111_1111111111111111_1111101000101010_0101000000001000"; -- -0.02279186062514782
	pesos_i(3216) := b"1111111111111111_1111111111111111_1111000001101011_0100001111010000"; -- -0.06086326763033867
	pesos_i(3217) := b"0000000000000000_0000000000000000_0000011111110010_1000001011100000"; -- 0.03104417771100998
	pesos_i(3218) := b"0000000000000000_0000000000000000_0100011010101101_0011011110000000"; -- 0.27608057856559753
	pesos_i(3219) := b"0000000000000000_0000000000000000_0001110000111011_0010010001000000"; -- 0.11027742922306061
	pesos_i(3220) := b"1111111111111111_1111111111111111_1110101111011110_0010111000000000"; -- -0.07864105701446533
	pesos_i(3221) := b"1111111111111111_1111111111111111_1110101011110010_0011010001000000"; -- -0.08224175870418549
	pesos_i(3222) := b"1111111111111111_1111111111111111_1111001111100111_1110000011010000"; -- -0.04724306985735893
	pesos_i(3223) := b"0000000000000000_0000000000000000_0001010111010110_0011000010100000"; -- 0.0852995291352272
	pesos_i(3224) := b"1111111111111111_1111111111111111_1101100010110111_1100111101000000"; -- -0.1534452885389328
	pesos_i(3225) := b"0000000000000000_0000000000000000_0001111100100110_1101000111100000"; -- 0.12168609350919724
	pesos_i(3226) := b"0000000000000000_0000000000000000_0000010000001000_0000011101111000"; -- 0.015747515484690666
	pesos_i(3227) := b"1111111111111111_1111111111111111_1111111100001000_1001101111001000"; -- -0.0037748944014310837
	pesos_i(3228) := b"0000000000000000_0000000000000000_0011110010000010_0101101010000000"; -- 0.23636403679847717
	pesos_i(3229) := b"0000000000000000_0000000000000000_0000110111010001_0111110111000000"; -- 0.053977832198143005
	pesos_i(3230) := b"0000000000000000_0000000000000000_0000110000001100_0000101111100000"; -- 0.04705881327390671
	pesos_i(3231) := b"0000000000000000_0000000000000000_0001110011100110_1010011000000000"; -- 0.11289441585540771
	pesos_i(3232) := b"1111111111111111_1111111111111111_1110000111010100_0001110100100000"; -- -0.11785715073347092
	pesos_i(3233) := b"0000000000000000_0000000000000000_0001011001010100_0000111101000000"; -- 0.08722014725208282
	pesos_i(3234) := b"1111111111111111_1111111111111111_1110110100010011_0111001100000000"; -- -0.07392197847366333
	pesos_i(3235) := b"1111111111111111_1111111111111111_1111101010110111_1101100000000000"; -- -0.020632266998291016
	pesos_i(3236) := b"0000000000000000_0000000000000000_0000101101101100_1010010001100000"; -- 0.044626496732234955
	pesos_i(3237) := b"1111111111111111_1111111111111111_1111010100000001_0011101101110000"; -- -0.04294994845986366
	pesos_i(3238) := b"1111111111111111_1111111111111111_1010111010101100_0101111100000000"; -- -0.31768232583999634
	pesos_i(3239) := b"0000000000000000_0000000000000000_0010111001000110_0110110111000000"; -- 0.1807621568441391
	pesos_i(3240) := b"0000000000000000_0000000000000000_0000011010100100_1000111001010000"; -- 0.025948423892259598
	pesos_i(3241) := b"0000000000000000_0000000000000000_0010111001010101_0010000100000000"; -- 0.1809864640235901
	pesos_i(3242) := b"0000000000000000_0000000000000000_0001001001010100_1010100011100000"; -- 0.07160430401563644
	pesos_i(3243) := b"1111111111111111_1111111111111111_1110000010111110_1111010001100000"; -- -0.12208626419305801
	pesos_i(3244) := b"0000000000000000_0000000000000000_0010010110101010_0010111110000000"; -- 0.14712807536125183
	pesos_i(3245) := b"1111111111111111_1111111111111111_1100100100011010_1000110110000000"; -- -0.21443858742713928
	pesos_i(3246) := b"0000000000000000_0000000000000000_0011000110111110_0010001001000000"; -- 0.19430746138095856
	pesos_i(3247) := b"0000000000000000_0000000000000000_0000010111001111_0000011001000000"; -- 0.022690191864967346
	pesos_i(3248) := b"1111111111111111_1111111111111111_1101110101001000_1101001001000000"; -- -0.13560758531093597
	pesos_i(3249) := b"1111111111111111_1111111111111111_1100101001011011_1010011101000000"; -- -0.20953898131847382
	pesos_i(3250) := b"1111111111111111_1111111111111111_1100000011101001_1000011010000000"; -- -0.2464366853237152
	pesos_i(3251) := b"0000000000000000_0000000000000000_0010000101100110_0111000101000000"; -- 0.1304693967103958
	pesos_i(3252) := b"0000000000000000_0000000000000000_0100010011011111_0101000010000000"; -- 0.2690325081348419
	pesos_i(3253) := b"1111111111111111_1111111111111111_1101101010000100_0111111001000000"; -- -0.1464158147573471
	pesos_i(3254) := b"1111111111111111_1111111111111111_1110110101110111_1100111001000000"; -- -0.07239066064357758
	pesos_i(3255) := b"1111111111111111_1111111111111111_1100100111101110_1110001111000000"; -- -0.2111985832452774
	pesos_i(3256) := b"1111111111111111_1111111111111111_1100110110100101_1100011100000000"; -- -0.1966891884803772
	pesos_i(3257) := b"0000000000000000_0000000000000000_0011010111111101_0100010001000000"; -- 0.21089579164981842
	pesos_i(3258) := b"0000000000000000_0000000000000000_0000000001001101_0100100100101010"; -- 0.001179287675768137
	pesos_i(3259) := b"0000000000000000_0000000000000000_0011001011001111_1111010101000000"; -- 0.19848568737506866
	pesos_i(3260) := b"0000000000000000_0000000000000000_0010000010000110_1000011111000000"; -- 0.12705276906490326
	pesos_i(3261) := b"0000000000000000_0000000000000000_0010101001101011_0110111000000000"; -- 0.1657017469406128
	pesos_i(3262) := b"1111111111111111_1111111111111111_1101100010011000_1111101111000000"; -- -0.1539156585931778
	pesos_i(3263) := b"1111111111111111_1111111111111111_1101110100010101_1000110011000000"; -- -0.13638992607593536
	pesos_i(3264) := b"0000000000000000_0000000000000000_0000101101000010_1010100111100000"; -- 0.04398595541715622
	pesos_i(3265) := b"0000000000000000_0000000000000000_0000000101010101_0010000111010000"; -- 0.005205262452363968
	pesos_i(3266) := b"1111111111111111_1111111111111111_1110110011111111_1111100011100000"; -- -0.07421917468309402
	pesos_i(3267) := b"1111111111111111_1111111111111111_1110000011101101_1011101000000000"; -- -0.12137258052825928
	pesos_i(3268) := b"0000000000000000_0000000000000000_0010101110100000_1100101011000000"; -- 0.1704222410917282
	pesos_i(3269) := b"1111111111111111_1111111111111111_1011111101010001_1010111010000000"; -- -0.2526598870754242
	pesos_i(3270) := b"1111111111111111_1111111111111111_1001001011010111_1111010000000000"; -- -0.4263923168182373
	pesos_i(3271) := b"0000000000000000_0000000000000000_0000110000111000_0001100010000000"; -- 0.047730952501297
	pesos_i(3272) := b"1111111111111111_1111111111111111_1001111101100000_1000000000000000"; -- -0.37743377685546875
	pesos_i(3273) := b"0000000000000000_0000000000000000_0001001101111100_0101110101000000"; -- 0.0761163979768753
	pesos_i(3274) := b"1111111111111111_1111111111111111_1110111111101101_1001011100100000"; -- -0.06278090924024582
	pesos_i(3275) := b"0000000000000000_0000000000000000_0001101001111011_1010110011100000"; -- 0.10344963520765305
	pesos_i(3276) := b"0000000000000000_0000000000000000_0011100111100010_0111101010000000"; -- 0.22611203789710999
	pesos_i(3277) := b"0000000000000000_0000000000000000_0011100100000100_0101111111000000"; -- 0.22272299230098724
	pesos_i(3278) := b"1111111111111111_1111111111111111_1100010011010001_1111111011000000"; -- -0.23117072880268097
	pesos_i(3279) := b"1111111111111111_1111111111111111_1000101000101010_0001001100000000"; -- -0.46029549837112427
	pesos_i(3280) := b"1111111111111111_1111111111111111_1101001101011011_0000001110000000"; -- -0.1743924915790558
	pesos_i(3281) := b"0000000000000000_0000000000000000_0010101111011000_1000101010000000"; -- 0.1712729036808014
	pesos_i(3282) := b"1111111111111111_1111111111111111_1110001100111001_1001001011000000"; -- -0.11240275204181671
	pesos_i(3283) := b"0000000000000000_0000000000000000_0000110000110110_1110110100110000"; -- 0.04771311208605766
	pesos_i(3284) := b"0000000000000000_0000000000000000_0011100100010010_0000110111000000"; -- 0.22293172776699066
	pesos_i(3285) := b"0000000000000000_0000000000000000_0001001101011010_0000000100100000"; -- 0.07559210807085037
	pesos_i(3286) := b"0000000000000000_0000000000000000_0001101010111110_0010010100100000"; -- 0.10446388274431229
	pesos_i(3287) := b"1111111111111111_1111111111111111_1111010110101000_1100110000010000"; -- -0.04039311036467552
	pesos_i(3288) := b"0000000000000000_0000000000000000_0011100000101101_0110101000000000"; -- 0.2194429636001587
	pesos_i(3289) := b"1111111111111111_1111111111111111_1110011100101111_0110011000100000"; -- -0.09693299978971481
	pesos_i(3290) := b"0000000000000000_0000000000000000_0001100101001001_0101100111100000"; -- 0.09877549856901169
	pesos_i(3291) := b"1111111111111111_1111111111111111_1001010110110010_1010101010000000"; -- -0.4152425229549408
	pesos_i(3292) := b"0000000000000000_0000000000000000_0000100101100100_0111111111100000"; -- 0.03668975085020065
	pesos_i(3293) := b"1111111111111111_1111111111111111_1111011101011101_1101001000110000"; -- -0.03372465446591377
	pesos_i(3294) := b"1111111111111111_1111111111111111_1111110011101001_1010001000010100"; -- -0.012060041539371014
	pesos_i(3295) := b"0000000000000000_0000000000000000_0000101001001001_1100101110010000"; -- 0.04018852487206459
	pesos_i(3296) := b"1111111111111111_1111111111111111_1101001001000001_0100101111000000"; -- -0.17869116365909576
	pesos_i(3297) := b"0000000000000000_0000000000000000_0000011110110011_1010001101000000"; -- 0.030084803700447083
	pesos_i(3298) := b"0000000000000000_0000000000000000_0001010000111100_0110100111000000"; -- 0.079046830534935
	pesos_i(3299) := b"1111111111111111_1111111111111111_1100000101101000_0001111000000000"; -- -0.24450504779815674
	pesos_i(3300) := b"0000000000000000_0000000000000000_0000110100111000_0010011100000000"; -- 0.05163806676864624
	pesos_i(3301) := b"0000000000000000_0000000000000000_0010000100101011_1011101110000000"; -- 0.12957355380058289
	pesos_i(3302) := b"1111111111111111_1111111111111111_1110110101011010_0011111111100000"; -- -0.07284165173768997
	pesos_i(3303) := b"1111111111111111_1111111111111111_0110111001110111_1001001000000000"; -- -0.5684880018234253
	pesos_i(3304) := b"0000000000000000_0000000000000000_0001001101100110_1110100100100000"; -- 0.07578904181718826
	pesos_i(3305) := b"0000000000000000_0000000000000000_0001011110111000_0111010000100000"; -- 0.09265828877687454
	pesos_i(3306) := b"1111111111111111_1111111111111111_1110111010100100_0001010011100000"; -- -0.06780881434679031
	pesos_i(3307) := b"1111111111111111_1111111111111111_1111101000001011_0000100001101000"; -- -0.023269152268767357
	pesos_i(3308) := b"1111111111111111_1111111111111111_1100110000011100_0110111100000000"; -- -0.20269113779067993
	pesos_i(3309) := b"1111111111111111_1111111111111111_1011001110101111_1011000000000000"; -- -0.29810047149658203
	pesos_i(3310) := b"0000000000000000_0000000000000000_0000010101111000_0011101100111000"; -- 0.021365834400057793
	pesos_i(3311) := b"1111111111111111_1111111111111111_1101001110110111_1110010010000000"; -- -0.17297527194023132
	pesos_i(3312) := b"1111111111111111_1111111111111111_1111110111010101_0001111001110000"; -- -0.008466813713312149
	pesos_i(3313) := b"1111111111111111_1111111111111111_0010110001110011_0101110000000000"; -- -0.8263647556304932
	pesos_i(3314) := b"1111111111111111_1111111111111111_1011110000111101_0101100010000000"; -- -0.2646889388561249
	pesos_i(3315) := b"1111111111111111_1111111111111111_1111110000011000_1101100101100100"; -- -0.015245831571519375
	pesos_i(3316) := b"1111111111111111_1111111111111111_1111110100000101_1001101001111100"; -- -0.011633248068392277
	pesos_i(3317) := b"0000000000000000_0000000000000000_0010101101111001_0111011110000000"; -- 0.16982218623161316
	pesos_i(3318) := b"1111111111111111_1111111111111111_1011100101011110_1000000010000000"; -- -0.27590176463127136
	pesos_i(3319) := b"0000000000000000_0000000000000000_0000110001100000_0001101000000000"; -- 0.04834139347076416
	pesos_i(3320) := b"1111111111111111_1111111111111111_1111111011011000_0001110010001000"; -- -0.004514900967478752
	pesos_i(3321) := b"1111111111111111_1111111111111111_1100000010110010_0101001101000000"; -- -0.24727897346019745
	pesos_i(3322) := b"1111111111111111_1111111111111111_1111101110010110_0000000110101000"; -- -0.01724233292043209
	pesos_i(3323) := b"1111111111111111_1111111111111111_1110011011010111_0000101110100000"; -- -0.09828116744756699
	pesos_i(3324) := b"0000000000000000_0000000000000000_0001011010011011_1010000010000000"; -- 0.08831217885017395
	pesos_i(3325) := b"1111111111111111_1111111111111111_1110011101101111_0111001000100000"; -- -0.09595572203397751
	pesos_i(3326) := b"0000000000000000_0000000000000000_0010111011011100_0111110101000000"; -- 0.18305189907550812
	pesos_i(3327) := b"1111111111111111_1111111111111111_1110100011111001_0110010001100000"; -- -0.08994457870721817
	pesos_i(3328) := b"1111111111111111_1111111111111111_1010110000100101_1100100000000000"; -- -0.3275485038757324
	pesos_i(3329) := b"1111111111111111_1111111111111111_1111111000010010_1111001100010000"; -- -0.007523354142904282
	pesos_i(3330) := b"1111111111111111_1111111111111111_1011000110111111_1001111110000000"; -- -0.3056698143482208
	pesos_i(3331) := b"0000000000000000_0000000000000000_0101000101100100_0111001010000000"; -- 0.3179389536380768
	pesos_i(3332) := b"1111111111111111_1111111111111111_1011101010110110_1001100110000000"; -- -0.270651251077652
	pesos_i(3333) := b"0000000000000000_0000000000000000_0100100000101101_1111011010000000"; -- 0.28195133805274963
	pesos_i(3334) := b"1111111111111111_1111111111111111_1101011010100110_0111110110000000"; -- -0.1615220606327057
	pesos_i(3335) := b"0000000000000000_0000000000000000_0001001100101010_0001001011000000"; -- 0.07486073672771454
	pesos_i(3336) := b"0000000000000000_0000000000000000_0100011101100111_0000101000000000"; -- 0.27891600131988525
	pesos_i(3337) := b"0000000000000000_0000000000000000_0010101101011001_1111100111000000"; -- 0.16934166848659515
	pesos_i(3338) := b"0000000000000000_0000000000000000_0010000101001010_1001100101000000"; -- 0.13004453480243683
	pesos_i(3339) := b"1111111111111111_1111111111111111_1011010011101111_1111100100000000"; -- -0.2932133078575134
	pesos_i(3340) := b"0000000000000000_0000000000000000_1000100011110110_0110101000000000"; -- 0.5350099802017212
	pesos_i(3341) := b"0000000000000000_0000000000000000_0001011010010110_0111010011000000"; -- 0.08823327720165253
	pesos_i(3342) := b"1111111111111111_1111111111111111_1101010101011101_1000010111000000"; -- -0.1665417104959488
	pesos_i(3343) := b"0000000000000000_0000000000000000_0011000100001101_0011010010000000"; -- 0.1916077435016632
	pesos_i(3344) := b"0000000000000000_0000000000000000_0001111111110000_1111110011000000"; -- 0.12477092444896698
	pesos_i(3345) := b"1111111111111111_1111111111111111_1101000001000101_1000010000000000"; -- -0.18643927574157715
	pesos_i(3346) := b"0000000000000000_0000000000000000_0001110110000100_0101010000100000"; -- 0.11530042439699173
	pesos_i(3347) := b"0000000000000000_0000000000000000_0001010101110001_1010100111000000"; -- 0.08376561105251312
	pesos_i(3348) := b"0000000000000000_0000000000000000_0001011010010100_0010011010100000"; -- 0.08819810301065445
	pesos_i(3349) := b"1111111111111111_1111111111111111_1100111110110101_1010011000000000"; -- -0.18863451480865479
	pesos_i(3350) := b"0000000000000000_0000000000000000_0011010000011110_0100010001000000"; -- 0.20358683168888092
	pesos_i(3351) := b"0000000000000000_0000000000000000_0101011101010101_1111011000000000"; -- 0.34115540981292725
	pesos_i(3352) := b"0000000000000000_0000000000000000_0100001001010010_0010001100000000"; -- 0.25906580686569214
	pesos_i(3353) := b"0000000000000000_0000000000000000_0110010101111101_0111001100000000"; -- 0.39644545316696167
	pesos_i(3354) := b"1111111111111111_1111111111111111_1001001111100110_1011000000000000"; -- -0.42226123809814453
	pesos_i(3355) := b"1111111111111111_1111111111111111_1111101001110011_1111110011010000"; -- -0.02166767045855522
	pesos_i(3356) := b"0000000000000000_0000000000000000_0110001100010000_0111111110000000"; -- 0.38697049021720886
	pesos_i(3357) := b"0000000000000000_0000000000000000_0011000110011010_0111001011000000"; -- 0.19376294314861298
	pesos_i(3358) := b"1111111111111111_1111111111111111_1110010001110010_1001010111100000"; -- -0.10762656480073929
	pesos_i(3359) := b"0000000000000000_0000000000000000_0101011000010010_0011111100000000"; -- 0.33621591329574585
	pesos_i(3360) := b"0000000000000000_0000000000000000_0001111011000001_1010010110000000"; -- 0.12014231085777283
	pesos_i(3361) := b"0000000000000000_0000000000000000_0000111011010111_0000010001010000"; -- 0.057968396693468094
	pesos_i(3362) := b"1111111111111111_1111111111111111_1111000110101000_1001000111010000"; -- -0.05602158233523369
	pesos_i(3363) := b"0000000000000000_0000000000000000_0010100011101101_0000001000000000"; -- 0.15986645221710205
	pesos_i(3364) := b"1111111111111111_1111111111111111_1100010010110001_0100100001000000"; -- -0.23166988790035248
	pesos_i(3365) := b"1111111111111111_1111111111111111_1101001010100011_0101100100000000"; -- -0.1771950125694275
	pesos_i(3366) := b"1111111111111111_1111111111111111_1100111110100101_0001001011000000"; -- -0.18888743221759796
	pesos_i(3367) := b"0000000000000000_0000000000000000_0111000000111101_0100100110000000"; -- 0.4384351670742035
	pesos_i(3368) := b"0000000000000000_0000000000000000_0000101001101111_0110111110110000"; -- 0.04076288267970085
	pesos_i(3369) := b"0000000000000000_0000000000000000_0000000101110010_0110011101001000"; -- 0.005651907995343208
	pesos_i(3370) := b"1111111111111111_1111111111111111_1111110011011011_0100000101101000"; -- -0.01227942667901516
	pesos_i(3371) := b"0000000000000000_0000000000000000_0010101010000111_0100011001000000"; -- 0.16612662374973297
	pesos_i(3372) := b"0000000000000000_0000000000000000_0000010000000111_0001101101111000"; -- 0.015733448788523674
	pesos_i(3373) := b"1111111111111111_1111111111111111_1111110100100011_0010111000011000"; -- -0.011181944981217384
	pesos_i(3374) := b"0000000000000000_0000000000000000_0101000000010110_0000000100000000"; -- 0.3128357529640198
	pesos_i(3375) := b"0000000000000000_0000000000000000_0000110010101000_1001111111110000"; -- 0.049448009580373764
	pesos_i(3376) := b"1111111111111111_1111111111111111_1100011011000000_0001010011000000"; -- -0.2236315757036209
	pesos_i(3377) := b"1111111111111111_1111111111111111_1001011100100000_0101011010000000"; -- -0.40966281294822693
	pesos_i(3378) := b"0000000000000000_0000000000000000_0011101101000110_1001000100000000"; -- 0.23154550790786743
	pesos_i(3379) := b"1111111111111111_1111111111111111_1111111101111010_0001101101101011"; -- -0.0020430434960871935
	pesos_i(3380) := b"0000000000000000_0000000000000000_0101101011101100_1101110000000000"; -- 0.3551766872406006
	pesos_i(3381) := b"0000000000000000_0000000000000000_0010111000101100_0100100101000000"; -- 0.1803632527589798
	pesos_i(3382) := b"1111111111111111_1111111111111111_1111010011111011_1101001101000000"; -- -0.0430324524641037
	pesos_i(3383) := b"1111111111111111_1111111111111111_1001100100111100_0011100110000000"; -- -0.4014247953891754
	pesos_i(3384) := b"0000000000000000_0000000000000000_0110000001110101_0001000000000000"; -- 0.3767862319946289
	pesos_i(3385) := b"1111111111111111_1111111111111111_1011111011100011_1101010010000000"; -- -0.25433608889579773
	pesos_i(3386) := b"0000000000000000_0000000000000000_0110010111000100_1101111100000000"; -- 0.3975352644920349
	pesos_i(3387) := b"1111111111111111_1111111111111111_1100011011011011_1111111110000000"; -- -0.2232055962085724
	pesos_i(3388) := b"1111111111111111_1111111111111111_1101100000001101_0010100011000000"; -- -0.1560492068529129
	pesos_i(3389) := b"0000000000000000_0000000000000000_0100011100111010_0101000010000000"; -- 0.2782335579395294
	pesos_i(3390) := b"1111111111111111_1111111111111111_1101010010110000_1010001110000000"; -- -0.16917970776557922
	pesos_i(3391) := b"0000000000000000_0000000000000000_0001111000110010_0010011100000000"; -- 0.11795276403427124
	pesos_i(3392) := b"0000000000000000_0000000000000000_0010011111101100_0100111101000000"; -- 0.15594954788684845
	pesos_i(3393) := b"1111111111111111_1111111111111111_1111010011011010_1110110000100000"; -- -0.04353450983762741
	pesos_i(3394) := b"0000000000000000_0000000000000000_0000000110110100_1111110000111000"; -- 0.006667865440249443
	pesos_i(3395) := b"1111111111111111_1111111111111111_1110011001011011_0001001100000000"; -- -0.10017281770706177
	pesos_i(3396) := b"1111111111111111_1111111111111111_1100111111000111_1100011000000000"; -- -0.18835794925689697
	pesos_i(3397) := b"1111111111111111_1111111111111111_1001001100011111_0001100100000000"; -- -0.4253067374229431
	pesos_i(3398) := b"1111111111111111_1111111111111111_1100111111010001_1001011010000000"; -- -0.1882081925868988
	pesos_i(3399) := b"0000000000000000_0000000000000000_0000101101000010_1111101100010000"; -- 0.04399079456925392
	pesos_i(3400) := b"0000000000000000_0000000000000000_0011001101111110_1011111000000000"; -- 0.20115268230438232
	pesos_i(3401) := b"0000000000000000_0000000000000000_0110001110000111_1110110010000000"; -- 0.3887927830219269
	pesos_i(3402) := b"0000000000000000_0000000000000000_0001111000101111_0011101111100000"; -- 0.11790823191404343
	pesos_i(3403) := b"1111111111111111_1111111111111111_1111100000101001_0110011100010000"; -- -0.030618246644735336
	pesos_i(3404) := b"0000000000000000_0000000000000000_0000101110101111_1110110100000000"; -- 0.04565316438674927
	pesos_i(3405) := b"1111111111111111_1111111111111111_1110001101010101_0000111001100000"; -- -0.11198339611291885
	pesos_i(3406) := b"1111111111111111_1111111111111111_1100010100110010_0010111101000000"; -- -0.22970299422740936
	pesos_i(3407) := b"1111111111111111_1111111111111111_1001001101110100_0010111000000000"; -- -0.42400848865509033
	pesos_i(3408) := b"0000000000000000_0000000000000000_0001110100001110_1010111000000000"; -- 0.11350524425506592
	pesos_i(3409) := b"0000000000000000_0000000000000000_0010010100011000_0001010000000000"; -- 0.1448986530303955
	pesos_i(3410) := b"0000000000000000_0000000000000000_0011001011110111_0110110010000000"; -- 0.19908788800239563
	pesos_i(3411) := b"0000000000000000_0000000000000000_0011100001101111_0011111011000000"; -- 0.22044746577739716
	pesos_i(3412) := b"0000000000000000_0000000000000000_0011001001000111_0100101011000000"; -- 0.19640032947063446
	pesos_i(3413) := b"0000000000000000_0000000000000000_0011000001011001_0011011011000000"; -- 0.18886129558086395
	pesos_i(3414) := b"0000000000000000_0000000000000000_0001011001110010_1110011011100000"; -- 0.08769076317548752
	pesos_i(3415) := b"0000000000000000_0000000000000000_0001010100100000_0001000000100000"; -- 0.082520492374897
	pesos_i(3416) := b"0000000000000000_0000000000000000_0011111101101111_0110000000000000"; -- 0.24779319763183594
	pesos_i(3417) := b"1111111111111111_1111111111111111_1111110011100001_0011000100000000"; -- -0.012188851833343506
	pesos_i(3418) := b"1111111111111111_1111111111111111_1110001001111011_1111000100100000"; -- -0.11529629677534103
	pesos_i(3419) := b"1111111111111111_1111111111111111_1101100000111001_0100110101000000"; -- -0.1553756445646286
	pesos_i(3420) := b"1111111111111111_1111111111111111_1110110110110101_0100100010100000"; -- -0.07145258039236069
	pesos_i(3421) := b"0000000000000000_0000000000000000_0100010010111000_1000110000000000"; -- 0.26844096183776855
	pesos_i(3422) := b"0000000000000000_0000000000000000_0011111011111111_0100110100000000"; -- 0.2460830807685852
	pesos_i(3423) := b"1111111111111111_1111111111111111_1101010110100000_0000011000000000"; -- -0.16552698612213135
	pesos_i(3424) := b"1111111111111111_1111111111111111_1010110010110001_1110001100000000"; -- -0.3254106640815735
	pesos_i(3425) := b"1111111111111111_1111111111111111_1110110101010110_1000010111100000"; -- -0.0728985145688057
	pesos_i(3426) := b"1111111111111111_1111111111111111_1101101100000011_1111101010000000"; -- -0.14447054266929626
	pesos_i(3427) := b"0000000000000000_0000000000000000_0001100111110011_0001011011000000"; -- 0.10136549174785614
	pesos_i(3428) := b"1111111111111111_1111111111111111_1111110111011011_0110011000110100"; -- -0.00837098341435194
	pesos_i(3429) := b"0000000000000000_0000000000000000_0000010011101111_1001101101000000"; -- 0.01928110420703888
	pesos_i(3430) := b"1111111111111111_1111111111111111_1110000101000110_1011010111000000"; -- -0.12001480162143707
	pesos_i(3431) := b"1111111111111111_1111111111111111_0101000101100001_0000101000000000"; -- -0.6821130514144897
	pesos_i(3432) := b"0000000000000000_0000000000000000_0100000111101001_0000011010000000"; -- 0.25746193528175354
	pesos_i(3433) := b"0000000000000000_0000000000000000_0000111000001010_1001011010000000"; -- 0.054849058389663696
	pesos_i(3434) := b"0000000000000000_0000000000000000_0001111000001001_0001001100100000"; -- 0.11732596904039383
	pesos_i(3435) := b"0000000000000000_0000000000000000_0000000000101001_1010100010100101"; -- 0.0006356623489409685
	pesos_i(3436) := b"1111111111111111_1111111111111111_1100011110001001_1010100110000000"; -- -0.22055569291114807
	pesos_i(3437) := b"0000000000000000_0000000000000000_0011010101111111_1001110101000000"; -- 0.20897848904132843
	pesos_i(3438) := b"1111111111111111_1111111111111111_1101011101111000_0110111101000000"; -- -0.15831856429576874
	pesos_i(3439) := b"1111111111111111_1111111111111111_1100101100111101_1011001101000000"; -- -0.2060897797346115
	pesos_i(3440) := b"1111111111111111_1111111111111111_1110000101011111_0101010001100000"; -- -0.11963913589715958
	pesos_i(3441) := b"1111111111111111_1111111111111111_0011101110101110_0110110100000000"; -- -0.7668697237968445
	pesos_i(3442) := b"1111111111111111_1111111111111111_1110111010110100_0110101110000000"; -- -0.06755951046943665
	pesos_i(3443) := b"1111111111111111_1111111111111111_1101001100110100_1100001011000000"; -- -0.17497618496418
	pesos_i(3444) := b"0000000000000000_0000000000000000_0011101011111100_0111111111000000"; -- 0.23041532933712006
	pesos_i(3445) := b"0000000000000000_0000000000000000_0100111000011100_0011010110000000"; -- 0.3051179349422455
	pesos_i(3446) := b"1111111111111111_1111111111111111_1100011010000100_0101000111000000"; -- -0.2245434671640396
	pesos_i(3447) := b"1111111111111111_1111111111111111_1100111001000001_1000111011000000"; -- -0.1943121701478958
	pesos_i(3448) := b"0000000000000000_0000000000000000_0001111011101110_0001101000000000"; -- 0.12082064151763916
	pesos_i(3449) := b"1111111111111111_1111111111111111_1110101011001110_1101100100000000"; -- -0.08278125524520874
	pesos_i(3450) := b"0000000000000000_0000000000000000_0100111000101110_1000000010000000"; -- 0.30539706349372864
	pesos_i(3451) := b"0000000000000000_0000000000000000_0110000110000101_1010100010000000"; -- 0.38094571232795715
	pesos_i(3452) := b"0000000000000000_0000000000000000_0011010000010110_1011010011000000"; -- 0.20347146689891815
	pesos_i(3453) := b"0000000000000000_0000000000000000_0000110100100010_1110000000110000"; -- 0.05131341144442558
	pesos_i(3454) := b"0000000000000000_0000000000000000_0001010011101010_0111000101100000"; -- 0.08170231431722641
	pesos_i(3455) := b"1111111111111111_1111111111111111_1110110111011000_0100100100000000"; -- -0.0709185004234314
	pesos_i(3456) := b"0000000000000000_0000000000000000_0001110011010001_0011010001000000"; -- 0.11256720125675201
	pesos_i(3457) := b"1111111111111111_1111111111111111_1111110101011100_0011001011100100"; -- -0.010311908088624477
	pesos_i(3458) := b"1111111111111111_1111111111111111_1100010101001000_0000111000000000"; -- -0.22936928272247314
	pesos_i(3459) := b"0000000000000000_0000000000000000_0101110011111110_0011100110000000"; -- 0.3632541596889496
	pesos_i(3460) := b"1111111111111111_1111111111111111_1011010001111011_1010101100000000"; -- -0.2949879765510559
	pesos_i(3461) := b"0000000000000000_0000000000000000_0011111110110101_1001010111000000"; -- 0.24886451661586761
	pesos_i(3462) := b"0000000000000000_0000000000000000_0100101010010000_1010011110000000"; -- 0.2912697494029999
	pesos_i(3463) := b"0000000000000000_0000000000000000_0001110001101110_1110011000000000"; -- 0.11106717586517334
	pesos_i(3464) := b"0000000000000000_0000000000000000_0000101011010011_0110101101000000"; -- 0.04228849709033966
	pesos_i(3465) := b"0000000000000000_0000000000000000_0110111000101011_0111000110000000"; -- 0.4303503930568695
	pesos_i(3466) := b"0000000000000000_0000000000000000_0010110001011010_1001000010000000"; -- 0.17325690388679504
	pesos_i(3467) := b"1111111111111111_1111111111111111_1010111111000111_1100010000000000"; -- -0.3133580684661865
	pesos_i(3468) := b"0000000000000000_0000000000000000_0100110100101010_0000011010000000"; -- 0.30142250657081604
	pesos_i(3469) := b"0000000000000000_0000000000000000_0001111101111010_0111101000100000"; -- 0.1229626014828682
	pesos_i(3470) := b"1111111111111111_1111111111111111_1111111110011010_0101111111001110"; -- -0.0015506859635934234
	pesos_i(3471) := b"0000000000000000_0000000000000000_0011010100011011_1001100000000000"; -- 0.20745229721069336
	pesos_i(3472) := b"1111111111111111_1111111111111111_1110010001101110_0010000110100000"; -- -0.10769452899694443
	pesos_i(3473) := b"0000000000000000_0000000000000000_0011011101001011_0000101100000000"; -- 0.21598881483078003
	pesos_i(3474) := b"1111111111111111_1111111111111111_1100100101111000_1101010000000000"; -- -0.21300005912780762
	pesos_i(3475) := b"1111111111111111_1111111111111111_1000010110110101_1110001100000000"; -- -0.4776933789253235
	pesos_i(3476) := b"0000000000000000_0000000000000000_0001010110110100_1101100101100000"; -- 0.08479078859090805
	pesos_i(3477) := b"1111111111111111_1111111111111111_1110001101101000_0011011110000000"; -- -0.11169102787971497
	pesos_i(3478) := b"0000000000000000_0000000000000000_0000011001011010_0110001101001000"; -- 0.024816708639264107
	pesos_i(3479) := b"0000000000000000_0000000000000000_0001101011010000_1011101010100000"; -- 0.10474745184183121
	pesos_i(3480) := b"0000000000000000_0000000000000000_0101000111110001_0110010010000000"; -- 0.3200896084308624
	pesos_i(3481) := b"0000000000000000_0000000000000000_0011001000110100_1011101101000000"; -- 0.1961171180009842
	pesos_i(3482) := b"0000000000000000_0000000000000000_0011010101101001_1100011100000000"; -- 0.2086452841758728
	pesos_i(3483) := b"1111111111111111_1111111111111111_1011111110010011_0100100100000000"; -- -0.2516588568687439
	pesos_i(3484) := b"0000000000000000_0000000000000000_1000101001101100_1101100000000000"; -- 0.5407233238220215
	pesos_i(3485) := b"0000000000000000_0000000000000000_0001100110110001_0011000000100000"; -- 0.10035992413759232
	pesos_i(3486) := b"0000000000000000_0000000000000000_0011100101111101_1100100101000000"; -- 0.22457559406757355
	pesos_i(3487) := b"0000000000000000_0000000000000000_0000010110101110_0010101001110000"; -- 0.022188808768987656
	pesos_i(3488) := b"0000000000000000_0000000000000000_1000010101110111_0010010000000000"; -- 0.5213491916656494
	pesos_i(3489) := b"1111111111111111_1111111111111111_1001110111010010_1001111000000000"; -- -0.3835049867630005
	pesos_i(3490) := b"0000000000000000_0000000000000000_0100011111011101_1000010110000000"; -- 0.28072389960289
	pesos_i(3491) := b"0000000000000000_0000000000000000_0011101110000111_1111110100000000"; -- 0.23254376649856567
	pesos_i(3492) := b"0000000000000000_0000000000000000_0111010001001010_1101111110000000"; -- 0.4542674720287323
	pesos_i(3493) := b"0000000000000000_0000000000000000_0010110110110001_1111010010000000"; -- 0.17849662899971008
	pesos_i(3494) := b"0000000000000000_0000000000000000_0111101100001110_0111100110000000"; -- 0.4806896150112152
	pesos_i(3495) := b"0000000000000000_0000000000000000_0010000110011011_0110100100000000"; -- 0.13127762079238892
	pesos_i(3496) := b"0000000000000000_0000000000000000_0100010100010101_1001101010000000"; -- 0.2698608934879303
	pesos_i(3497) := b"1111111111111111_1111111111111111_1101011001100110_0010100001000000"; -- -0.1625037044286728
	pesos_i(3498) := b"0000000000000000_0000000000000000_0100001010111110_0111100100000000"; -- 0.2607188820838928
	pesos_i(3499) := b"0000000000000000_0000000000000000_0101000110010010_1010111010000000"; -- 0.3186444342136383
	pesos_i(3500) := b"0000000000000000_0000000000000000_0000000010000100_1010110100000111"; -- 0.002024473389610648
	pesos_i(3501) := b"1111111111111111_1111111111111111_1100011001110111_0110101000000000"; -- -0.2247403860092163
	pesos_i(3502) := b"1111111111111111_1111111111111111_1110101111100111_0001101111000000"; -- -0.07850481569766998
	pesos_i(3503) := b"0000000000000000_0000000000000000_0010001001010001_1010101100000000"; -- 0.1340586543083191
	pesos_i(3504) := b"0000000000000000_0000000000000000_0011101100010001_1000001011000000"; -- 0.23073594272136688
	pesos_i(3505) := b"1111111111111111_1111111111111111_0110001111010010_0001011100000000"; -- -0.6100755333900452
	pesos_i(3506) := b"0000000000000000_0000000000000000_0110110010011010_1101001110000000"; -- 0.424237459897995
	pesos_i(3507) := b"1111111111111111_1111111111111111_1101110001101011_0111110010000000"; -- -0.13898488879203796
	pesos_i(3508) := b"0000000000000000_0000000000000000_0011110000010010_0111110101000000"; -- 0.23465712368488312
	pesos_i(3509) := b"0000000000000000_0000000000000000_0101111000000100_1110111000000000"; -- 0.36726272106170654
	pesos_i(3510) := b"0000000000000000_0000000000000000_0000110010111110_0011101001110000"; -- 0.04977765306830406
	pesos_i(3511) := b"1111111111111111_1111111111111111_1111010010100111_1011110001110000"; -- -0.04431555047631264
	pesos_i(3512) := b"0000000000000000_0000000000000000_0110001010010001_1001100010000000"; -- 0.38503411412239075
	pesos_i(3513) := b"1111111111111111_1111111111111111_1101111100011010_0001110101000000"; -- -0.12850777804851532
	pesos_i(3514) := b"0000000000000000_0000000000000000_0001010110110011_0011101110000000"; -- 0.08476611971855164
	pesos_i(3515) := b"0000000000000000_0000000000000000_0000110101111100_0010101011010000"; -- 0.052675891667604446
	pesos_i(3516) := b"1111111111111111_1111111111111111_1111100100111001_1010101101111000"; -- -0.02646377868950367
	pesos_i(3517) := b"1111111111111111_1111111111111111_1110111101100100_0100010011000000"; -- -0.06487627327442169
	pesos_i(3518) := b"1111111111111111_1111111111111111_1101011111010101_1001000101000000"; -- -0.15689747035503387
	pesos_i(3519) := b"1111111111111111_1111111111111111_1101000011111100_0000011000000000"; -- -0.18365442752838135
	pesos_i(3520) := b"0000000000000000_0000000000000000_0001001111010110_0111111101000000"; -- 0.07749171555042267
	pesos_i(3521) := b"0000000000000000_0000000000000000_0001110010001100_0001010010100000"; -- 0.11151245981454849
	pesos_i(3522) := b"0000000000000000_0000000000000000_0010010111101000_0100001111000000"; -- 0.14807532727718353
	pesos_i(3523) := b"0000000000000000_0000000000000000_0010001100011001_1111111001000000"; -- 0.13711537420749664
	pesos_i(3524) := b"0000000000000000_0000000000000000_0000010011010101_1001000111010000"; -- 0.01888381317257881
	pesos_i(3525) := b"1111111111111111_1111111111111111_0111101100000101_0101001100000000"; -- -0.5194500088691711
	pesos_i(3526) := b"0000000000000000_0000000000000000_1000110101010011_1111011000000000"; -- 0.5520623922348022
	pesos_i(3527) := b"1111111111111111_1111111111111111_1110100001110100_1111001001100000"; -- -0.09196553379297256
	pesos_i(3528) := b"0000000000000000_0000000000000000_0011010110000101_0100011111000000"; -- 0.20906494557857513
	pesos_i(3529) := b"1111111111111111_1111111111111111_1100101111010010_0001011010000000"; -- -0.20382556319236755
	pesos_i(3530) := b"0000000000000000_0000000000000000_0101101001100111_1111011100000000"; -- 0.353148877620697
	pesos_i(3531) := b"0000000000000000_0000000000000000_0110010000110100_1010111000000000"; -- 0.3914288282394409
	pesos_i(3532) := b"0000000000000000_0000000000000000_0001000010011010_0001000111000000"; -- 0.06485091149806976
	pesos_i(3533) := b"1111111111111111_1111111111111111_1110010101100000_0000001010000000"; -- -0.10400375723838806
	pesos_i(3534) := b"0000000000000000_0000000000000000_1010100111001111_0010111000000000"; -- 0.6633175611495972
	pesos_i(3535) := b"0000000000000000_0000000000000000_1011011001101100_0101111000000000"; -- 0.7125910520553589
	pesos_i(3536) := b"1111111111111111_1111111111111111_1100001000010011_0101111101000000"; -- -0.24189190566539764
	pesos_i(3537) := b"1111111111111111_1111111111111111_1111011000110110_1101100101000000"; -- -0.038225576281547546
	pesos_i(3538) := b"0000000000000000_0000000000000000_0000001001110101_0100111011010000"; -- 0.00960247591137886
	pesos_i(3539) := b"1111111111111111_1111111111111111_1111101001101110_0111100000100000"; -- -0.021751873195171356
	pesos_i(3540) := b"0000000000000000_0000000000000000_0010000001010000_1111100110000000"; -- 0.12623557448387146
	pesos_i(3541) := b"0000000000000000_0000000000000000_0101001011100010_0100000110000000"; -- 0.3237648904323578
	pesos_i(3542) := b"1111111111111111_1111111111111111_1111101011100110_0101011110100000"; -- -0.019922755658626556
	pesos_i(3543) := b"1111111111111111_1111111111111111_0111011011010101_1100100100000000"; -- -0.5358003973960876
	pesos_i(3544) := b"0000000000000000_0000000000000000_0000011100100111_0011110100101000"; -- 0.027942487969994545
	pesos_i(3545) := b"0000000000000000_0000000000000000_0100100101010011_1011111000000000"; -- 0.2864340543746948
	pesos_i(3546) := b"1111111111111111_1111111111111111_1111011011001101_1011010011000000"; -- -0.03592367470264435
	pesos_i(3547) := b"1111111111111111_1111111111111111_1011101110011011_1011001110000000"; -- -0.2671554386615753
	pesos_i(3548) := b"1111111111111111_1111111111111111_1001000000001100_0010011110000000"; -- -0.43731454014778137
	pesos_i(3549) := b"0000000000000000_0000000000000000_0000001101101110_1001000100010000"; -- 0.01340586319565773
	pesos_i(3550) := b"0000000000000000_0000000000000000_0001010010101011_0011101001000000"; -- 0.08073772490024567
	pesos_i(3551) := b"1111111111111111_1111111111111111_1100001111101000_0010100001000000"; -- -0.2347388118505478
	pesos_i(3552) := b"1111111111111111_1111111111111111_1100010000001101_1110000110000000"; -- -0.23416319489479065
	pesos_i(3553) := b"0000000000000000_0000000000000000_0000010000101001_0100010101000000"; -- 0.016254737973213196
	pesos_i(3554) := b"1111111111111111_1111111111111111_1101000110110010_0011000101000000"; -- -0.1808747500181198
	pesos_i(3555) := b"0000000000000000_0000000000000000_1000111110011011_1101111000000000"; -- 0.5609720945358276
	pesos_i(3556) := b"0000000000000000_0000000000000000_0001111100000010_1101110011100000"; -- 0.12113743275403976
	pesos_i(3557) := b"1111111111111111_1111111111111111_1000000000010100_1101000010000000"; -- -0.49968239665031433
	pesos_i(3558) := b"0000000000000000_0000000000000000_0100101011011101_1111101000000000"; -- 0.29244959354400635
	pesos_i(3559) := b"1111111111111111_1111111111111110_1001100010101001_1001010000000000"; -- -1.4036624431610107
	pesos_i(3560) := b"0000000000000000_0000000000000000_0101100011001101_0100110100000000"; -- 0.3468826413154602
	pesos_i(3561) := b"1111111111111111_1111111111111111_1111001101100011_1000101111000000"; -- -0.04926230013370514
	pesos_i(3562) := b"1111111111111111_1111111111111111_1011010010111100_1011011100000000"; -- -0.2939954400062561
	pesos_i(3563) := b"0000000000000000_0000000000000000_0000101010010110_0110110111100000"; -- 0.041357867419719696
	pesos_i(3564) := b"0000000000000000_0000000000000000_0101010010001011_0001101100000000"; -- 0.33024758100509644
	pesos_i(3565) := b"0000000000000000_0000000000000000_0110000111110110_1100000100000000"; -- 0.38267141580581665
	pesos_i(3566) := b"1111111111111111_1111111111111111_1001111000010011_0000011100000000"; -- -0.3825221657752991
	pesos_i(3567) := b"1111111111111111_1111111111111111_0110100000011000_0001111000000000"; -- -0.5933820009231567
	pesos_i(3568) := b"0000000000000000_0000000000000000_0011001010111001_1001001010000000"; -- 0.1981441080570221
	pesos_i(3569) := b"1111111111111111_1111111111111111_1000111101111101_0110010110000000"; -- -0.4394928514957428
	pesos_i(3570) := b"1111111111111111_1111111111111111_1111111111000110_0101011101111101"; -- -0.0008797951159067452
	pesos_i(3571) := b"1111111111111111_1111111111111111_1010010010111010_1011101010000000"; -- -0.3565257489681244
	pesos_i(3572) := b"0000000000000000_0000000000000000_0011001001110101_1000101001000000"; -- 0.1971060186624527
	pesos_i(3573) := b"1111111111111111_1111111111111111_1011001000000001_0111100100000000"; -- -0.3046650290489197
	pesos_i(3574) := b"1111111111111111_1111111111111111_0110011100001000_0110000100000000"; -- -0.5975283980369568
	pesos_i(3575) := b"0000000000000000_0000000000000000_0000010100010101_1100100110111000"; -- 0.019863707944750786
	pesos_i(3576) := b"0000000000000000_0000000000000000_0100001011101001_1011110110000000"; -- 0.26137909293174744
	pesos_i(3577) := b"1111111111111111_1111111111111111_1111000111111000_0010010001000000"; -- -0.05480740964412689
	pesos_i(3578) := b"0000000000000000_0000000000000000_0101010100001111_0001011010000000"; -- 0.33226147294044495
	pesos_i(3579) := b"1111111111111111_1111111111111111_1111010110010011_0010100111100000"; -- -0.04072321206331253
	pesos_i(3580) := b"0000000000000000_0000000000000000_0110011010110100_0011001010000000"; -- 0.40118709206581116
	pesos_i(3581) := b"0000000000000000_0000000000000000_0010101111100111_1100100001000000"; -- 0.17150546610355377
	pesos_i(3582) := b"1111111111111111_1111111111111111_1110010111011111_1101100101100000"; -- -0.10205308347940445
	pesos_i(3583) := b"1111111111111111_1111111111111111_1000100110001100_1101011010000000"; -- -0.4626947343349457
	pesos_i(3584) := b"0000000000000000_0000000000000000_0011101111011010_1111111100000000"; -- 0.23381036520004272
	pesos_i(3585) := b"0000000000000000_0000000000000000_0001010110110011_1000101101100000"; -- 0.08477088063955307
	pesos_i(3586) := b"1111111111111111_1111111111111111_1001101111000101_1011000100000000"; -- -0.39151471853256226
	pesos_i(3587) := b"1111111111111111_1111111111111111_1000111010110000_0101100000000000"; -- -0.44262170791625977
	pesos_i(3588) := b"0000000000000000_0000000000000000_0110111111110100_1010000100000000"; -- 0.43732649087905884
	pesos_i(3589) := b"0000000000000000_0000000000000000_0110110111000101_1101100110000000"; -- 0.42880019545555115
	pesos_i(3590) := b"1111111111111111_1111111111111111_1100110001010011_0000110010000000"; -- -0.2018577754497528
	pesos_i(3591) := b"0000000000000000_0000000000000000_0100010111101100_0101001100000000"; -- 0.27313727140426636
	pesos_i(3592) := b"0000000000000000_0000000000000000_0111111001101010_0100100000000000"; -- 0.49380922317504883
	pesos_i(3593) := b"1111111111111111_1111111111111111_1100010101000011_0100000010000000"; -- -0.2294425666332245
	pesos_i(3594) := b"0000000000000000_0000000000000000_0001100110001011_0101010101000000"; -- 0.0997823029756546
	pesos_i(3595) := b"0000000000000000_0000000000000000_0110110011110111_1100011010000000"; -- 0.4256557524204254
	pesos_i(3596) := b"1111111111111111_1111111111111111_1100000010010000_0011000101000000"; -- -0.2477997988462448
	pesos_i(3597) := b"1111111111111111_1111111111111111_1110111100000100_1111111011100000"; -- -0.06633002310991287
	pesos_i(3598) := b"1111111111111111_1111111111111111_0111101010000100_0001011000000000"; -- -0.5214220285415649
	pesos_i(3599) := b"0000000000000000_0000000000000000_0101011001011011_1101101000000000"; -- 0.33733904361724854
	pesos_i(3600) := b"0000000000000000_0000000000000000_0011111110110011_1010001110000000"; -- 0.24883481860160828
	pesos_i(3601) := b"1111111111111111_1111111111111111_1111101010111011_1100110101001000"; -- -0.020571870729327202
	pesos_i(3602) := b"1111111111111111_1111111111111111_1110111011110100_1010011001000000"; -- -0.06657944619655609
	pesos_i(3603) := b"1111111111111111_1111111111111111_1110000000100100_1001000011000000"; -- -0.12444205582141876
	pesos_i(3604) := b"1111111111111111_1111111111111111_1010110100010111_0101001000000000"; -- -0.3238629102706909
	pesos_i(3605) := b"0000000000000000_0000000000000000_0111010110011011_0010001100000000"; -- 0.45939844846725464
	pesos_i(3606) := b"1111111111111111_1111111111111111_1000011010010110_0100100010000000"; -- -0.4742693603038788
	pesos_i(3607) := b"0000000000000000_0000000000000000_1000110010001101_1010010100000000"; -- 0.5490363240242004
	pesos_i(3608) := b"1111111111111111_1111111111111111_1100010100100100_0110110101000000"; -- -0.2299129217863083
	pesos_i(3609) := b"1111111111111111_1111111111111111_1110000001011000_1001110110000000"; -- -0.12364783883094788
	pesos_i(3610) := b"0000000000000000_0000000000000000_0111100110011110_0110010000000000"; -- 0.47507309913635254
	pesos_i(3611) := b"0000000000000000_0000000000000000_0010111010010001_0000001110000000"; -- 0.1819002330303192
	pesos_i(3612) := b"0000000000000000_0000000000000000_1000000000010111_0001111000000000"; -- 0.5003527402877808
	pesos_i(3613) := b"1111111111111111_1111111111111111_0111101010011011_1101111000000000"; -- -0.5210591554641724
	pesos_i(3614) := b"0000000000000000_0000000000000000_0100011011001110_1010100010000000"; -- 0.27659085392951965
	pesos_i(3615) := b"0000000000000000_0000000000000000_0000110100001101_0001011010010000"; -- 0.050980959087610245
	pesos_i(3616) := b"0000000000000000_0000000000000000_0101010010010001_0001000010000000"; -- 0.3303385078907013
	pesos_i(3617) := b"1111111111111111_1111111111111111_0100110100000001_0011101000000000"; -- -0.6992000341415405
	pesos_i(3618) := b"1111111111111111_1111111111111111_1101010101010101_0011000110000000"; -- -0.16666880249977112
	pesos_i(3619) := b"1111111111111111_1111111111111111_1011111111111001_1100111000000000"; -- -0.25009453296661377
	pesos_i(3620) := b"0000000000000000_0000000000000000_0110001100001011_1111000010000000"; -- 0.386900931596756
	pesos_i(3621) := b"0000000000000000_0000000000000000_0101101110001010_1011100100000000"; -- 0.35758548974990845
	pesos_i(3622) := b"0000000000000000_0000000000000000_0110001011110110_0111100100000000"; -- 0.3865733742713928
	pesos_i(3623) := b"1111111111111111_1111111111111111_1011000100001000_1001001010000000"; -- -0.3084629476070404
	pesos_i(3624) := b"1111111111111111_1111111111111111_1011001100101000_0100001000000000"; -- -0.3001669645309448
	pesos_i(3625) := b"0000000000000000_0000000000000000_0100111001111001_1110111110000000"; -- 0.3065480887889862
	pesos_i(3626) := b"0000000000000000_0000000000000000_0001001000101100_1111110100000000"; -- 0.07099896669387817
	pesos_i(3627) := b"0000000000000000_0000000000000000_0100001111111010_1100110110000000"; -- 0.26554569602012634
	pesos_i(3628) := b"0000000000000000_0000000000000000_0111111111111000_0010101010000000"; -- 0.49988046288490295
	pesos_i(3629) := b"1111111111111111_1111111111111111_1000010100110100_1101010100000000"; -- -0.47966259717941284
	pesos_i(3630) := b"0000000000000000_0000000000000000_0001111001000110_0111111001100000"; -- 0.11826314777135849
	pesos_i(3631) := b"1111111111111111_1111111111111111_1001011001110100_0010011110000000"; -- -0.41229012608528137
	pesos_i(3632) := b"0000000000000000_0000000000000000_0011101000111110_0100000100000000"; -- 0.2275124192237854
	pesos_i(3633) := b"0000000000000000_0000000000000000_0110001010101111_0100010000000000"; -- 0.3854868412017822
	pesos_i(3634) := b"0000000000000000_0000000000000000_0110010111010000_0000000100000000"; -- 0.3977051377296448
	pesos_i(3635) := b"0000000000000000_0000000000000000_0011100110000101_0100111001000000"; -- 0.22469033300876617
	pesos_i(3636) := b"1111111111111111_1111111111111111_1100011010101001_1010011100000000"; -- -0.22397381067276
	pesos_i(3637) := b"0000000000000000_0000000000000000_0101010000010000_1100100010000000"; -- 0.32838109135627747
	pesos_i(3638) := b"1111111111111111_1111111111111111_1110001110001000_0001110001000000"; -- -0.1112043708562851
	pesos_i(3639) := b"1111111111111111_1111111111111111_1110100011000101_1001101110100000"; -- -0.09073474258184433
	pesos_i(3640) := b"0000000000000000_0000000000000000_0100110111010101_0001101100000000"; -- 0.30403298139572144
	pesos_i(3641) := b"0000000000000000_0000000000000000_0101101001110100_0011000100000000"; -- 0.353335440158844
	pesos_i(3642) := b"0000000000000000_0000000000000000_0100000000001101_1001111100000000"; -- 0.2502078413963318
	pesos_i(3643) := b"0000000000000000_0000000000000000_0011100110001010_1111001001000000"; -- 0.22477640211582184
	pesos_i(3644) := b"0000000000000000_0000000000000000_0101100111101100_1010011100000000"; -- 0.3512672781944275
	pesos_i(3645) := b"1111111111111111_1111111111111111_1001101010011000_0011010010000000"; -- -0.3961150348186493
	pesos_i(3646) := b"1111111111111111_1111111111111111_1111001110000010_0011001011110000"; -- -0.048794571310281754
	pesos_i(3647) := b"1111111111111111_1111111111111111_1101111100000010_0100010101000000"; -- -0.1288716048002243
	pesos_i(3648) := b"1111111111111111_1111111111111111_0110011000110100_1101011100000000"; -- -0.6007562279701233
	pesos_i(3649) := b"0000000000000000_0000000000000000_0101101110011010_1111000110000000"; -- 0.35783299803733826
	pesos_i(3650) := b"0000000000000000_0000000000000000_0110001110111001_0101111000000000"; -- 0.3895472288131714
	pesos_i(3651) := b"1111111111111111_1111111111111111_0110100011111000_1010011100000000"; -- -0.5899558663368225
	pesos_i(3652) := b"0000000000000000_0000000000000000_0111000001010101_1011001110000000"; -- 0.4388076961040497
	pesos_i(3653) := b"0000000000000000_0000000000000000_0101100111000000_1101101110000000"; -- 0.3505990207195282
	pesos_i(3654) := b"0000000000000000_0000000000000000_0001010011010010_0111101100000000"; -- 0.08133667707443237
	pesos_i(3655) := b"1111111111111111_1111111111111111_1011111100101111_0111101010000000"; -- -0.2531817853450775
	pesos_i(3656) := b"1111111111111111_1111111111111111_1011110000111100_1001010010000000"; -- -0.26470062136650085
	pesos_i(3657) := b"1111111111111111_1111111111111111_0110011001111001_0010111100000000"; -- -0.5997133851051331
	pesos_i(3658) := b"0000000000000000_0000000000000000_0101010111111101_1110001110000000"; -- 0.3359052836894989
	pesos_i(3659) := b"0000000000000000_0000000000000000_0111100111011001_0110011110000000"; -- 0.47597357630729675
	pesos_i(3660) := b"0000000000000000_0000000000000000_0000011111101100_1101101100111000"; -- 0.030957890674471855
	pesos_i(3661) := b"1111111111111111_1111111111111111_1101101100001110_0101011011000000"; -- -0.14431245625019073
	pesos_i(3662) := b"0000000000000000_0000000000000000_0010011001100100_1010000001000000"; -- 0.14997293055057526
	pesos_i(3663) := b"0000000000000000_0000000000000000_0111010000101101_1111110100000000"; -- 0.4538267254829407
	pesos_i(3664) := b"1111111111111111_1111111111111111_1100001000011110_1010000110000000"; -- -0.24172011017799377
	pesos_i(3665) := b"0000000000000000_0000000000000000_0110011010100000_1101011100000000"; -- 0.4008917212486267
	pesos_i(3666) := b"0000000000000000_0000000000000000_0000110101011101_1101010010100000"; -- 0.05221299082040787
	pesos_i(3667) := b"1111111111111111_1111111111111111_0110000111101010_0110001000000000"; -- -0.617517352104187
	pesos_i(3668) := b"1111111111111111_1111111111111111_1100101110111110_1010001001000000"; -- -0.2041224092245102
	pesos_i(3669) := b"0000000000000000_0000000000000000_0000100111111101_1110111100100000"; -- 0.039030976593494415
	pesos_i(3670) := b"1111111111111111_1111111111111111_1100000110110100_1111101100000000"; -- -0.24333220720291138
	pesos_i(3671) := b"1111111111111111_1111111111111111_1110000110101111_1100011000000000"; -- -0.11841166019439697
	pesos_i(3672) := b"1111111111111111_1111111111111111_1111010010101100_1100101010000000"; -- -0.04423841834068298
	pesos_i(3673) := b"1111111111111111_1111111111111111_1110111100100011_0000101111000000"; -- -0.06587149202823639
	pesos_i(3674) := b"0000000000000000_0000000000000000_0001001100011100_1111000100100000"; -- 0.07466036826372147
	pesos_i(3675) := b"1111111111111111_1111111111111111_1001101000010101_1000101000000000"; -- -0.3981088399887085
	pesos_i(3676) := b"0000000000000000_0000000000000000_0001101111011100_1011100010000000"; -- 0.10883668065071106
	pesos_i(3677) := b"1111111111111111_1111111111111111_1100111100100100_0101010111000000"; -- -0.1908518224954605
	pesos_i(3678) := b"0000000000000000_0000000000000000_0110101011001011_1111100100000000"; -- 0.4171748757362366
	pesos_i(3679) := b"0000000000000000_0000000000000000_0001010100100000_0000111100100000"; -- 0.08252043277025223
	pesos_i(3680) := b"0000000000000000_0000000000000000_0010010011011011_0100110001000000"; -- 0.14397121965885162
	pesos_i(3681) := b"0000000000000000_0000000000000000_0001001111011110_0010000111100000"; -- 0.07760822027921677
	pesos_i(3682) := b"1111111111111111_1111111111111111_1110001101100110_1100111010100000"; -- -0.11171253770589828
	pesos_i(3683) := b"0000000000000000_0000000000000000_0101000110010110_1101110000000000"; -- 0.3187081813812256
	pesos_i(3684) := b"0000000000000000_0000000000000000_0001101000101110_1001011101100000"; -- 0.10227342694997787
	pesos_i(3685) := b"1111111111111111_1111111111111111_0100111101000110_0010011000000000"; -- -0.6903358697891235
	pesos_i(3686) := b"0000000000000000_0000000000000000_0011001011001001_0010011101000000"; -- 0.19838185608386993
	pesos_i(3687) := b"0000000000000000_0000000000000000_0011011000111001_1111010001000000"; -- 0.2118218094110489
	pesos_i(3688) := b"1111111111111111_1111111111111111_1110011101001111_1101001000000000"; -- -0.09643828868865967
	pesos_i(3689) := b"0000000000000000_0000000000000000_0011000100001000_1001000011000000"; -- 0.19153694808483124
	pesos_i(3690) := b"1111111111111111_1111111111111111_1001110010111010_0001011000000000"; -- -0.38778555393218994
	pesos_i(3691) := b"1111111111111111_1111111111111111_1001100001110101_0000101000000000"; -- -0.40446412563323975
	pesos_i(3692) := b"1111111111111111_1111111111111111_1101001001010010_1001100001000000"; -- -0.17842720448970795
	pesos_i(3693) := b"1111111111111111_1111111111111111_1111010100000111_1011111110000000"; -- -0.04285052418708801
	pesos_i(3694) := b"1111111111111111_1111111111111111_1100001000010000_0010101101000000"; -- -0.24194078147411346
	pesos_i(3695) := b"1111111111111111_1111111111111111_1111011010111001_1100000101110000"; -- -0.03622809424996376
	pesos_i(3696) := b"0000000000000000_0000000000000000_0010000010001000_1010001001000000"; -- 0.1270848661661148
	pesos_i(3697) := b"0000000000000000_0000000000000000_0111110000101000_0111110110000000"; -- 0.4849928319454193
	pesos_i(3698) := b"0000000000000000_0000000000000000_0000100000111011_1100010100110000"; -- 0.03216202184557915
	pesos_i(3699) := b"0000000000000000_0000000000000000_0001110000101110_0111111110100000"; -- 0.11008451133966446
	pesos_i(3700) := b"0000000000000000_0000000000000000_0010100111000101_0010011001000000"; -- 0.16316451132297516
	pesos_i(3701) := b"1111111111111111_1111111111111111_1101111110001100_0001001000000000"; -- -0.12676894664764404
	pesos_i(3702) := b"1111111111111111_1111111111111111_1000100101001100_0001110000000000"; -- -0.4636824131011963
	pesos_i(3703) := b"0000000000000000_0000000000000000_0110011001101110_0011010000000000"; -- 0.4001190662384033
	pesos_i(3704) := b"0000000000000000_0000000000000000_0000110111000111_0001100111000000"; -- 0.053819283843040466
	pesos_i(3705) := b"1111111111111111_1111111111111111_1111111010000000_1001100100001000"; -- -0.005850253626704216
	pesos_i(3706) := b"0000000000000000_0000000000000000_0100010010010100_0000001010000000"; -- 0.26788344979286194
	pesos_i(3707) := b"0000000000000000_0000000000000000_0110000100010100_1011101110000000"; -- 0.3792226016521454
	pesos_i(3708) := b"1111111111111111_1111111111111111_1001010000111100_1000110000000000"; -- -0.42095112800598145
	pesos_i(3709) := b"0000000000000000_0000000000000000_0100001101010101_0010010010000000"; -- 0.2630179226398468
	pesos_i(3710) := b"1111111111111111_1111111111111111_1111101000011011_1001000010000000"; -- -0.023016899824142456
	pesos_i(3711) := b"1111111111111111_1111111111111111_1111011000010110_0100000101110000"; -- -0.03872290626168251
	pesos_i(3712) := b"1111111111111111_1111111111111111_1100110001011010_0011011111000000"; -- -0.20174838602542877
	pesos_i(3713) := b"1111111111111111_1111111111111111_1011011001100000_0101000000000000"; -- -0.28759288787841797
	pesos_i(3714) := b"0000000000000000_0000000000000000_0000101101110010_1101100011000000"; -- 0.044721171259880066
	pesos_i(3715) := b"0000000000000000_0000000000000000_0010111111010101_1110100010000000"; -- 0.18685773015022278
	pesos_i(3716) := b"0000000000000000_0000000000000000_0011000001111011_0001111111000000"; -- 0.18937872350215912
	pesos_i(3717) := b"1111111111111111_1111111111111111_1111111011000101_1010001001111010"; -- -0.004796834196895361
	pesos_i(3718) := b"0000000000000000_0000000000000000_0000111010111110_1101110100110000"; -- 0.05759985372424126
	pesos_i(3719) := b"1111111111111111_1111111111111111_1111110111100111_1001001101100000"; -- -0.008185185492038727
	pesos_i(3720) := b"0000000000000000_0000000000000000_0001111101011101_1011111001100000"; -- 0.12252416461706161
	pesos_i(3721) := b"1111111111111111_1111111111111111_1101101100000111_1001111001000000"; -- -0.1444150060415268
	pesos_i(3722) := b"1111111111111111_1111111111111111_1101000110100110_0111101110000000"; -- -0.18105342984199524
	pesos_i(3723) := b"0000000000000000_0000000000000000_0000011000100001_1100000110100000"; -- 0.023952580988407135
	pesos_i(3724) := b"0000000000000000_0000000000000000_0000110011000100_0110010100100000"; -- 0.04987175017595291
	pesos_i(3725) := b"0000000000000000_0000000000000000_0011001011000010_1100111000000000"; -- 0.19828498363494873
	pesos_i(3726) := b"1111111111111111_1111111111111111_1101100011011011_0000010110000000"; -- -0.15290799736976624
	pesos_i(3727) := b"0000000000000000_0000000000000000_0110111100011000_1011100000000000"; -- 0.43397092819213867
	pesos_i(3728) := b"0000000000000000_0000000000000000_0001110100111001_1011001101000000"; -- 0.11416168510913849
	pesos_i(3729) := b"1111111111111111_1111111111111111_1110001001001100_0101000111000000"; -- -0.11602295935153961
	pesos_i(3730) := b"1111111111111111_1111111111111111_1111110010010001_0110101010001000"; -- -0.013406125828623772
	pesos_i(3731) := b"1111111111111111_1111111111111111_1111101100000010_0001100000111000"; -- -0.019499288871884346
	pesos_i(3732) := b"1111111111111111_1111111111111111_1111110011110100_0100011011101100"; -- -0.01189762819558382
	pesos_i(3733) := b"0000000000000000_0000000000000000_0001110110111010_1111111100000000"; -- 0.11613458395004272
	pesos_i(3734) := b"1111111111111111_1111111111111111_1100101011000100_0011001111000000"; -- -0.20794369280338287
	pesos_i(3735) := b"0000000000000000_0000000000000000_0011011000100011_1100100000000000"; -- 0.21148347854614258
	pesos_i(3736) := b"1111111111111111_1111111111111111_1100011101111111_1010100011000000"; -- -0.22070832550525665
	pesos_i(3737) := b"0000000000000000_0000000000000000_0101110111000110_0111111110000000"; -- 0.36631008982658386
	pesos_i(3738) := b"1111111111111111_1111111111111111_1100100010100011_0000101111000000"; -- -0.2162621170282364
	pesos_i(3739) := b"0000000000000000_0000000000000000_0010010100001100_0011100001000000"; -- 0.14471770823001862
	pesos_i(3740) := b"0000000000000000_0000000000000000_0110101111101111_1000001010000000"; -- 0.4216233789920807
	pesos_i(3741) := b"1111111111111111_1111111111111111_1111111101000110_0111010001011011"; -- -0.002831199439242482
	pesos_i(3742) := b"1111111111111111_1111111111111111_1110000110111010_1011000011000000"; -- -0.11824508011341095
	pesos_i(3743) := b"0000000000000000_0000000000000000_0100111110001010_1101110110000000"; -- 0.31071266531944275
	pesos_i(3744) := b"0000000000000000_0000000000000000_0010110100100101_1011000001000000"; -- 0.17635633051395416
	pesos_i(3745) := b"1111111111111111_1111111111111111_1110001000011111_1111001001000000"; -- -0.11670003831386566
	pesos_i(3746) := b"1111111111111111_1111111111111111_1101100011001000_0110101101000000"; -- -0.15319184958934784
	pesos_i(3747) := b"1111111111111111_1111111111111111_1110010000010001_0111010011000000"; -- -0.10910864174365997
	pesos_i(3748) := b"1111111111111111_1111111111111111_1011000111000111_1111110010000000"; -- -0.3055422008037567
	pesos_i(3749) := b"1111111111111111_1111111111111111_1111101110101001_0110111001010000"; -- -0.016945939511060715
	pesos_i(3750) := b"1111111111111111_1111111111111111_1110010011001001_0101100001000000"; -- -0.10630272328853607
	pesos_i(3751) := b"0000000000000000_0000000000000000_0000010000100100_1010110100110000"; -- 0.016184639185667038
	pesos_i(3752) := b"1111111111111111_1111111111111111_0101011011111110_0000010100000000"; -- -0.6601864695549011
	pesos_i(3753) := b"1111111111111111_1111111111111111_1111110101010011_0101010001010000"; -- -0.010447245091199875
	pesos_i(3754) := b"1111111111111111_1111111111111111_1101110101000010_1010011010000000"; -- -0.1357017457485199
	pesos_i(3755) := b"0000000000000000_0000000000000000_0010001111000011_0000101111000000"; -- 0.1396949142217636
	pesos_i(3756) := b"1111111111111111_1111111111111111_1100101100111011_1010001011000000"; -- -0.2061212807893753
	pesos_i(3757) := b"1111111111111111_1111111111111111_1110010001010100_0011101111100000"; -- -0.10808969289064407
	pesos_i(3758) := b"0000000000000000_0000000000000000_0011111010101111_1000011010000000"; -- 0.2448658049106598
	pesos_i(3759) := b"1111111111111111_1111111111111111_1110010110111000_0010111001000000"; -- -0.10265837609767914
	pesos_i(3760) := b"1111111111111111_1111111111111111_1101100010101100_0100010111000000"; -- -0.15362133085727692
	pesos_i(3761) := b"1111111111111111_1111111111111111_1010000110001010_0000001110000000"; -- -0.3689878284931183
	pesos_i(3762) := b"0000000000000000_0000000000000000_0011001110111111_1101000001000000"; -- 0.20214559137821198
	pesos_i(3763) := b"0000000000000000_0000000000000000_0110101111111001_1101001110000000"; -- 0.4217807948589325
	pesos_i(3764) := b"0000000000000000_0000000000000000_0100100100010011_0100011100000000"; -- 0.28545039892196655
	pesos_i(3765) := b"0000000000000000_0000000000000000_0010100000100110_1011101010000000"; -- 0.1568409502506256
	pesos_i(3766) := b"1111111111111111_1111111111111111_1101010101000010_0100010001000000"; -- -0.16695760190486908
	pesos_i(3767) := b"0000000000000000_0000000000000000_0010000010111100_1111111010000000"; -- 0.12788382172584534
	pesos_i(3768) := b"1111111111111111_1111111111111111_1101010100101001_0010101001000000"; -- -0.16734062135219574
	pesos_i(3769) := b"1111111111111111_1111111111111111_1101010100101111_0100111100000000"; -- -0.16724687814712524
	pesos_i(3770) := b"0000000000000000_0000000000000000_0111011100100101_0111010000000000"; -- 0.46541523933410645
	pesos_i(3771) := b"1111111111111111_1111111111111111_1111101001001011_0010011110110000"; -- -0.022290725260972977
	pesos_i(3772) := b"1111111111111111_1111111111111111_1101100001110011_1000111000000000"; -- -0.1544867753982544
	pesos_i(3773) := b"1111111111111111_1111111111111111_1110110011001100_1110110011100000"; -- -0.07499808818101883
	pesos_i(3774) := b"0000000000000000_0000000000000000_0010010000101111_1010111010000000"; -- 0.1413525640964508
	pesos_i(3775) := b"0000000000000000_0000000000000000_0100001100001000_0000100000000000"; -- 0.2618412971496582
	pesos_i(3776) := b"1111111111111111_1111111111111111_0011101110110110_0110111000000000"; -- -0.7667475938796997
	pesos_i(3777) := b"1111111111111111_1111111111111111_1010011100001110_0101100110000000"; -- -0.3474372923374176
	pesos_i(3778) := b"1111111111111111_1111111111111111_1101110101001100_1011011100000000"; -- -0.1355481743812561
	pesos_i(3779) := b"1111111111111111_1111111111111111_1100100110011100_0001001000000000"; -- -0.21246230602264404
	pesos_i(3780) := b"1111111111111111_1111111111111111_1101100100000011_0010000001000000"; -- -0.1522960513830185
	pesos_i(3781) := b"1111111111111111_1111111111111111_1100110010000010_1000100011000000"; -- -0.20113320648670197
	pesos_i(3782) := b"1111111111111111_1111111111111111_1110100110010100_0100011101100000"; -- -0.08758119493722916
	pesos_i(3783) := b"0000000000000000_0000000000000000_0111000000000101_0101001000000000"; -- 0.4375811815261841
	pesos_i(3784) := b"0000000000000000_0000000000000000_0000011010000000_0100110011010000"; -- 0.02539520338177681
	pesos_i(3785) := b"0000000000000000_0000000000000000_0000001011101000_1001101010000100"; -- 0.011361748911440372
	pesos_i(3786) := b"0000000000000000_0000000000000000_0011010001000101_0010010010000000"; -- 0.2041800320148468
	pesos_i(3787) := b"1111111111111111_1111111111111111_1011101001100011_0000111010000000"; -- -0.27192601561546326
	pesos_i(3788) := b"1111111111111111_1111111111111111_1110011110101100_0101101100000000"; -- -0.09502631425857544
	pesos_i(3789) := b"0000000000000000_0000000000000000_1000100111011100_1100100100000000"; -- 0.5385251641273499
	pesos_i(3790) := b"1111111111111111_1111111111111111_1111001000011100_1100011110110000"; -- -0.054248351603746414
	pesos_i(3791) := b"1111111111111111_1111111111111111_1101111001101011_0000011001000000"; -- -0.13117943704128265
	pesos_i(3792) := b"0000000000000000_0000000000000000_0110111111101110_1001000000000000"; -- 0.43723392486572266
	pesos_i(3793) := b"0000000000000000_0000000000000000_0100001111011000_1000010010000000"; -- 0.26502254605293274
	pesos_i(3794) := b"0000000000000000_0000000000000000_0001111101100101_0101100110100000"; -- 0.1226402297616005
	pesos_i(3795) := b"1111111111111111_1111111111111111_1111111110100100_1100100011110010"; -- -0.0013918312033638358
	pesos_i(3796) := b"0000000000000000_0000000000000000_0010011100001011_1100011010000000"; -- 0.15252342820167542
	pesos_i(3797) := b"0000000000000000_0000000000000000_0001011010101011_1011001111000000"; -- 0.08855746686458588
	pesos_i(3798) := b"0000000000000000_0000000000000000_0100011101011001_1110011110000000"; -- 0.278715580701828
	pesos_i(3799) := b"0000000000000000_0000000000000000_0001001110110001_0010001011100000"; -- 0.07692163437604904
	pesos_i(3800) := b"0000000000000000_0000000000000000_0010100110111111_1101101100000000"; -- 0.1630837321281433
	pesos_i(3801) := b"0000000000000000_0000000000000000_0000111110101111_0100100011100000"; -- 0.06126838177442551
	pesos_i(3802) := b"0000000000000000_0000000000000000_1000010110010000_0110101100000000"; -- 0.521734893321991
	pesos_i(3803) := b"0000000000000000_0000000000000000_0010110111000100_1100101101000000"; -- 0.1787840873003006
	pesos_i(3804) := b"1111111111111111_1111111111111111_1110011010100000_1110110100000000"; -- -0.09910696744918823
	pesos_i(3805) := b"0000000000000000_0000000000000000_0101011100100011_1111110010000000"; -- 0.3403928577899933
	pesos_i(3806) := b"0000000000000000_0000000000000000_0010111100010000_1100110110000000"; -- 0.18385013937950134
	pesos_i(3807) := b"0000000000000000_0000000000000000_0001101111010011_0010011001000000"; -- 0.10869063436985016
	pesos_i(3808) := b"0000000000000000_0000000000000000_0000111010101110_1000011100000000"; -- 0.05735057592391968
	pesos_i(3809) := b"1111111111111111_1111111111111111_1101001101111110_0100000010000000"; -- -0.173854798078537
	pesos_i(3810) := b"0000000000000000_0000000000000000_0101101110010001_0101101100000000"; -- 0.35768669843673706
	pesos_i(3811) := b"1111111111111111_1111111111111111_1001101001100000_1101101110000000"; -- -0.3969595730304718
	pesos_i(3812) := b"0000000000000000_0000000000000000_0011111000001110_1011000111000000"; -- 0.24241171777248383
	pesos_i(3813) := b"1111111111111111_1111111111111111_1011100000110100_0000011010000000"; -- -0.28045615553855896
	pesos_i(3814) := b"1111111111111111_1111111111111111_1101110011001100_1001101010000000"; -- -0.1375029981136322
	pesos_i(3815) := b"0000000000000000_0000000000000000_0110000010111101_0110110010000000"; -- 0.37789037823677063
	pesos_i(3816) := b"0000000000000000_0000000000000000_0011100110100010_0111010000000000"; -- 0.22513508796691895
	pesos_i(3817) := b"1111111111111111_1111111111111111_0000001001111001_0001010000000000"; -- -0.990339994430542
	pesos_i(3818) := b"1111111111111111_1111111111111111_1101011111010101_1011010111000000"; -- -0.15689529478549957
	pesos_i(3819) := b"1111111111111111_1111111111111111_1110101011101111_0001001110000000"; -- -0.08228948712348938
	pesos_i(3820) := b"1111111111111111_1111111111111111_1001001110010010_0001011110000000"; -- -0.4235520660877228
	pesos_i(3821) := b"1111111111111111_1111111111111111_1101111100000010_0010100110000000"; -- -0.12887325882911682
	pesos_i(3822) := b"1111111111111111_1111111111111111_1111111110000100_1000101001011100"; -- -0.0018838430987671018
	pesos_i(3823) := b"0000000000000000_0000000000000000_0011000000100110_1100110101000000"; -- 0.18809206783771515
	pesos_i(3824) := b"1111111111111111_1111111111111111_1101000001010010_1000111110000000"; -- -0.18624022603034973
	pesos_i(3825) := b"1111111111111111_1111111111111111_1101101100101000_1011110100000000"; -- -0.14390963315963745
	pesos_i(3826) := b"1111111111111111_1111111111111111_1101100000010001_0011011000000000"; -- -0.15598738193511963
	pesos_i(3827) := b"0000000000000000_0000000000000000_0101110111001101_1001000010000000"; -- 0.36641791462898254
	pesos_i(3828) := b"1111111111111111_1111111111111111_1101011111110001_0001110100000000"; -- -0.156477153301239
	pesos_i(3829) := b"0000000000000000_0000000000000000_0001110100110011_0010001110000000"; -- 0.11406156420707703
	pesos_i(3830) := b"0000000000000000_0000000000000000_0011110000101100_1000110010000000"; -- 0.23505476117134094
	pesos_i(3831) := b"1111111111111111_1111111111111111_1111101010111101_1101001101010000"; -- -0.0205409936606884
	pesos_i(3832) := b"0000000000000000_0000000000000000_0000110001011000_0110111011000000"; -- 0.048224374651908875
	pesos_i(3833) := b"1111111111111111_1111111111111111_1111010101100011_0010111010100000"; -- -0.04145535081624985
	pesos_i(3834) := b"0000000000000000_0000000000000000_0000100111110111_1010010001000000"; -- 0.03893496096134186
	pesos_i(3835) := b"0000000000000000_0000000000000000_0010101000010000_0000010100000000"; -- 0.16430693864822388
	pesos_i(3836) := b"1111111111111111_1111111111111111_1101001111110110_1000101110000000"; -- -0.17201927304267883
	pesos_i(3837) := b"0000000000000000_0000000000000000_0100001000100110_1001111110000000"; -- 0.2584018409252167
	pesos_i(3838) := b"0000000000000000_0000000000000000_0010000000011100_1111001110000000"; -- 0.1254417598247528
	pesos_i(3839) := b"0000000000000000_0000000000000000_0100110100011100_1111011100000000"; -- 0.3012232184410095
	pesos_i(3840) := b"0000000000000000_0000000000000000_0000111010111001_0010111010010000"; -- 0.057513151317834854
	pesos_i(3841) := b"1111111111111111_1111111111111111_1011110100011111_0110101110000000"; -- -0.26123932003974915
	pesos_i(3842) := b"1111111111111111_1111111111111111_1110000111100101_1001010111000000"; -- -0.11759056150913239
	pesos_i(3843) := b"0000000000000000_0000000000000000_0001000110111010_0111001010100000"; -- 0.06925121694803238
	pesos_i(3844) := b"0000000000000000_0000000000000000_0001010100000000_1000101011000000"; -- 0.08203952014446259
	pesos_i(3845) := b"0000000000000000_0000000000000000_0011100100110000_1100101001000000"; -- 0.22340072691440582
	pesos_i(3846) := b"1111111111111111_1111111111111111_1100100000010011_0110000101000000"; -- -0.2184542864561081
	pesos_i(3847) := b"0000000000000000_0000000000000000_0011011100100110_1100011001000000"; -- 0.21543540060520172
	pesos_i(3848) := b"0000000000000000_0000000000000000_0001001001100001_1110101010100000"; -- 0.07180658727884293
	pesos_i(3849) := b"0000000000000000_0000000000000000_0001010011001000_1110111011100000"; -- 0.08119099587202072
	pesos_i(3850) := b"1111111111111111_1111111111111111_0101010111110111_1000010000000000"; -- -0.6641919612884521
	pesos_i(3851) := b"0000000000000000_0000000000000000_0001101100100100_0001101011100000"; -- 0.10601966828107834
	pesos_i(3852) := b"0000000000000000_0000000000000000_0001100111011000_1000001101100000"; -- 0.10095997899770737
	pesos_i(3853) := b"0000000000000000_0000000000000000_0001000010000010_1101011110000000"; -- 0.0644964873790741
	pesos_i(3854) := b"0000000000000000_0000000000000000_0100001001010001_0101101100000000"; -- 0.25905388593673706
	pesos_i(3855) := b"0000000000000000_0000000000000000_0010011011110101_1111001011000000"; -- 0.15219037234783173
	pesos_i(3856) := b"0000000000000000_0000000000000000_0011000111101000_0011000000000000"; -- 0.19494915008544922
	pesos_i(3857) := b"0000000000000000_0000000000000000_0001010000101111_0010101011000000"; -- 0.07884471118450165
	pesos_i(3858) := b"0000000000000000_0000000000000000_0010101111001110_0111111101000000"; -- 0.17111964523792267
	pesos_i(3859) := b"0000000000000000_0000000000000000_0100000111110010_1010100010000000"; -- 0.25760892033576965
	pesos_i(3860) := b"0000000000000000_0000000000000000_0010100111001110_1101000100000000"; -- 0.16331201791763306
	pesos_i(3861) := b"1111111111111111_1111111111111111_1111011100001010_0100110100100000"; -- -0.0349990651011467
	pesos_i(3862) := b"1111111111111111_1111111111111111_1110010111101011_0011100111100000"; -- -0.10187948495149612
	pesos_i(3863) := b"0000000000000000_0000000000000000_0000011011111001_0110110111110000"; -- 0.027243491262197495
	pesos_i(3864) := b"1111111111111111_1111111111111111_1110011111111110_0000100100100000"; -- -0.09377997368574142
	pesos_i(3865) := b"0000000000000000_0000000000000000_0100001000101100_1111110110000000"; -- 0.25849899649620056
	pesos_i(3866) := b"1111111111111111_1111111111111111_1011101001000101_1110000100000000"; -- -0.27237123250961304
	pesos_i(3867) := b"1111111111111111_1111111111111111_1110110010100111_0001011110000000"; -- -0.07557538151741028
	pesos_i(3868) := b"0000000000000000_0000000000000000_0111100111000010_0010111110000000"; -- 0.47561928629875183
	pesos_i(3869) := b"0000000000000000_0000000000000000_0101001001001110_0111001110000000"; -- 0.32150956988334656
	pesos_i(3870) := b"1111111111111111_1111111111111111_1111100110111010_0000100111110000"; -- -0.024505022913217545
	pesos_i(3871) := b"0000000000000000_0000000000000000_0110011111111111_0110010110000000"; -- 0.4062407910823822
	pesos_i(3872) := b"0000000000000000_0000000000000000_0010101001010001_0000001111000000"; -- 0.1652986854314804
	pesos_i(3873) := b"1111111111111111_1111111111111111_1100110100111101_1101111010000000"; -- -0.19827470183372498
	pesos_i(3874) := b"1111111111111111_1111111111111111_1111011011100101_0000010111000000"; -- -0.03556789457798004
	pesos_i(3875) := b"0000000000000000_0000000000000000_0001100000010111_0001010011100000"; -- 0.09410219639539719
	pesos_i(3876) := b"1111111111111111_1111111111111111_1101100000100100_0110111100000000"; -- -0.15569406747817993
	pesos_i(3877) := b"1111111111111111_1111111111111111_1110110010000011_1100110110100000"; -- -0.07611384242773056
	pesos_i(3878) := b"0000000000000000_0000000000000000_0000000000010000_1001111111011111"; -- 0.00025366965564899147
	pesos_i(3879) := b"1111111111111111_1111111111111111_1110011111000111_0111010101000000"; -- -0.09461276233196259
	pesos_i(3880) := b"1111111111111111_1111111111111110_1111000111101010_0100000000000000"; -- -1.0550193786621094
	pesos_i(3881) := b"0000000000000000_0000000000000000_0001011100000110_1111110001100000"; -- 0.08995034545660019
	pesos_i(3882) := b"0000000000000000_0000000000000000_0001101100101100_0100011110100000"; -- 0.10614440590143204
	pesos_i(3883) := b"0000000000000000_0000000000000000_0000111010101010_0101111011100000"; -- 0.057287149131298065
	pesos_i(3884) := b"1111111111111111_1111111111111111_1010010110111000_0110010000000000"; -- -0.35265517234802246
	pesos_i(3885) := b"0000000000000000_0000000000000000_0011100101111110_1011110111000000"; -- 0.22459016740322113
	pesos_i(3886) := b"0000000000000000_0000000000000000_0100001111110010_1000111010000000"; -- 0.2654198706150055
	pesos_i(3887) := b"1111111111111111_1111111111111111_1100011000011000_1011100011000000"; -- -0.22618527710437775
	pesos_i(3888) := b"0000000000000000_0000000000000000_0001001001001010_1101111100000000"; -- 0.07145494222640991
	pesos_i(3889) := b"0000000000000000_0000000000000000_0000110111100110_1100010110010000"; -- 0.05430254712700844
	pesos_i(3890) := b"1111111111111111_1111111111111111_1110110010000000_1101110000000000"; -- -0.07615876197814941
	pesos_i(3891) := b"0000000000000000_0000000000000000_0001101000110110_1110101000000000"; -- 0.10240042209625244
	pesos_i(3892) := b"0000000000000000_0000000000000000_0000011010010000_1010100101101000"; -- 0.02564486302435398
	pesos_i(3893) := b"0000000000000000_0000000000000000_0001111101011110_1111010110100000"; -- 0.12254271656274796
	pesos_i(3894) := b"0000000000000000_0000000000000000_0010000101101101_0010101100000000"; -- 0.13057202100753784
	pesos_i(3895) := b"1111111111111111_1111111111111111_1011110011110111_1101010000000000"; -- -0.2618434429168701
	pesos_i(3896) := b"1111111111111111_1111111111111111_1011111010011011_0110100100000000"; -- -0.2554411292076111
	pesos_i(3897) := b"1111111111111111_1111111111111111_1011111100100100_0000010110000000"; -- -0.25335660576820374
	pesos_i(3898) := b"0000000000000000_0000000000000000_0011010011001100_0101011001000000"; -- 0.20624293386936188
	pesos_i(3899) := b"1111111111111111_1111111111111111_1110001101000111_0101001000000000"; -- -0.11219298839569092
	pesos_i(3900) := b"0000000000000000_0000000000000000_0001000101100011_0100011000100000"; -- 0.06792104989290237
	pesos_i(3901) := b"0000000000000000_0000000000000000_0101111101100111_0101101000000000"; -- 0.3726707696914673
	pesos_i(3902) := b"1111111111111111_1111111111111111_1011101110000010_1110011010000000"; -- -0.2675338685512543
	pesos_i(3903) := b"0000000000000000_0000000000000000_0001110110111100_0011010011000000"; -- 0.1161530464887619
	pesos_i(3904) := b"1111111111111111_1111111111111111_0100100011011000_1111000000000000"; -- -0.7154397964477539
	pesos_i(3905) := b"1111111111111111_1111111111111111_1010111011000100_1111110000000000"; -- -0.3173067569732666
	pesos_i(3906) := b"1111111111111111_1111111111111111_1100001101101000_0000110101000000"; -- -0.23669354617595673
	pesos_i(3907) := b"0000000000000000_0000000000000000_0010011000100001_1110010110000000"; -- 0.14895471930503845
	pesos_i(3908) := b"1111111111111111_1111111111111111_1001011101000111_1100010000000000"; -- -0.4090611934661865
	pesos_i(3909) := b"0000000000000000_0000000000000000_0001100111000100_1111000110000000"; -- 0.10066136717796326
	pesos_i(3910) := b"1111111111111111_1111111111111111_1110111101000110_0011100001000000"; -- -0.06533478200435638
	pesos_i(3911) := b"0000000000000000_0000000000000000_0100000011110100_0010011100000000"; -- 0.25372546911239624
	pesos_i(3912) := b"0000000000000000_0000000000000000_0001001111000101_0011000000000000"; -- 0.07722759246826172
	pesos_i(3913) := b"1111111111111111_1111111111111111_1011010100001111_0100101110000000"; -- -0.29273536801338196
	pesos_i(3914) := b"1111111111111111_1111111111111111_1111000011110110_0001001010000000"; -- -0.058745235204696655
	pesos_i(3915) := b"0000000000000000_0000000000000000_0001001000000100_0101001101000000"; -- 0.07037849724292755
	pesos_i(3916) := b"0000000000000000_0000000000000000_0000101110101011_1000110111100000"; -- 0.04558645933866501
	pesos_i(3917) := b"0000000000000000_0000000000000000_0010001011011101_1110011111000000"; -- 0.1361985057592392
	pesos_i(3918) := b"0000000000000000_0000000000000000_0000000110110001_1000000110111000"; -- 0.006614787504076958
	pesos_i(3919) := b"1111111111111111_1111111111111111_1101111011101101_0110110001000000"; -- -0.12918971478939056
	pesos_i(3920) := b"1111111111111111_1111111111111111_1011100000100100_1011000000000000"; -- -0.28069019317626953
	pesos_i(3921) := b"1111111111111111_1111111111111111_1011100111000011_0001110010000000"; -- -0.2743665874004364
	pesos_i(3922) := b"0000000000000000_0000000000000000_0010011000101110_0111010001000000"; -- 0.14914633333683014
	pesos_i(3923) := b"0000000000000000_0000000000000000_0000000110010111_1111101000111110"; -- 0.006225242745131254
	pesos_i(3924) := b"1111111111111111_1111111111111111_1111110001110100_0010100001101100"; -- -0.01385257113724947
	pesos_i(3925) := b"1111111111111111_1111111111111111_1110010110101101_1110111111000000"; -- -0.1028146892786026
	pesos_i(3926) := b"1111111111111111_1111111111111111_1110111100000001_0100011100100000"; -- -0.06638675183057785
	pesos_i(3927) := b"1111111111111111_1111111111111111_1110011110110010_0111111000000000"; -- -0.0949326753616333
	pesos_i(3928) := b"1111111111111111_1111111111111111_1111001111111110_0110010010100000"; -- -0.046899519860744476
	pesos_i(3929) := b"0000000000000000_0000000000000000_0010010110011110_1011001110000000"; -- 0.14695283770561218
	pesos_i(3930) := b"1111111111111111_1111111111111111_1111011000111010_1000001011110000"; -- -0.03816968575119972
	pesos_i(3931) := b"1111111111111111_1111111111111111_1011111000011011_0001000110000000"; -- -0.25739946961402893
	pesos_i(3932) := b"1111111111111111_1111111111111111_1010001001110100_0001011100000000"; -- -0.36541610956192017
	pesos_i(3933) := b"0000000000000000_0000000000000000_0011010011000111_0001001100000000"; -- 0.20616263151168823
	pesos_i(3934) := b"0000000000000000_0000000000000000_0001000101100101_1100111011100000"; -- 0.06795971840620041
	pesos_i(3935) := b"1111111111111111_1111111111111111_1111101101100101_1111101101011000"; -- -0.017975131049752235
	pesos_i(3936) := b"0000000000000000_0000000000000000_0000100000001101_1110011100010000"; -- 0.031462136656045914
	pesos_i(3937) := b"1111111111111111_1111111111111111_1101011011000011_1000011010000000"; -- -0.1610790193080902
	pesos_i(3938) := b"0000000000000000_0000000000000000_0100010100110110_1010001100000000"; -- 0.2703649401664734
	pesos_i(3939) := b"1111111111111111_1111111111111111_0110001111001110_1111110000000000"; -- -0.6101229190826416
	pesos_i(3940) := b"0000000000000000_0000000000000000_0010010110100011_0101111010000000"; -- 0.14702406525611877
	pesos_i(3941) := b"0000000000000000_0000000000000000_0011010000100101_0001000000000000"; -- 0.2036905288696289
	pesos_i(3942) := b"1111111111111111_1111111111111111_1110010010011011_0010101110100000"; -- -0.10700728744268417
	pesos_i(3943) := b"0000000000000000_0000000000000000_0000010011101011_1111000111101000"; -- 0.019225234165787697
	pesos_i(3944) := b"1111111111111111_1111111111111111_1101010001100101_1001101010000000"; -- -0.1703246533870697
	pesos_i(3945) := b"1111111111111111_1111111111111110_1110001101000011_0001110000000000"; -- -1.1122572422027588
	pesos_i(3946) := b"1111111111111111_1111111111111111_1011110100001010_1000111000000000"; -- -0.2615576982498169
	pesos_i(3947) := b"0000000000000000_0000000000000000_0000101001000101_0101100011010000"; -- 0.040120650082826614
	pesos_i(3948) := b"1111111111111111_1111111111111111_1111101001101010_0111111101101000"; -- -0.021812474355101585
	pesos_i(3949) := b"1111111111111111_1111111111111111_0110011001001010_1001100100000000"; -- -0.6004242300987244
	pesos_i(3950) := b"0000000000000000_0000000000000000_0001000101011001_1110101001000000"; -- 0.06777824461460114
	pesos_i(3951) := b"1111111111111111_1111111111111111_1011001000011101_0111101110000000"; -- -0.30423763394355774
	pesos_i(3952) := b"0000000000000000_0000000000000000_0010011011001100_1100110001000000"; -- 0.15156246721744537
	pesos_i(3953) := b"1111111111111111_1111111111111111_1100011100010110_0010111000000000"; -- -0.22231781482696533
	pesos_i(3954) := b"1111111111111111_1111111111111111_1110001111011110_0011000010100000"; -- -0.1098909005522728
	pesos_i(3955) := b"1111111111111111_1111111111111111_1100100101101010_0010100100000000"; -- -0.2132238745689392
	pesos_i(3956) := b"0000000000000000_0000000000000000_0000010101111011_0111100110110000"; -- 0.021415334194898605
	pesos_i(3957) := b"0000000000000000_0000000000000000_0001111101110110_1011111111000000"; -- 0.12290571630001068
	pesos_i(3958) := b"1111111111111111_1111111111111111_1010111000000100_1000111010000000"; -- -0.3202429711818695
	pesos_i(3959) := b"1111111111111111_1111111111111111_0111000110011111_0110100000000000"; -- -0.5561614036560059
	pesos_i(3960) := b"0000000000000000_0000000000000000_0000000100010010_0100101101101110"; -- 0.004185404162853956
	pesos_i(3961) := b"0000000000000000_0000000000000000_0000010110111101_0111100010001000"; -- 0.022422345355153084
	pesos_i(3962) := b"0000000000000000_0000000000000000_0001000100011100_0000010010000000"; -- 0.06683376431465149
	pesos_i(3963) := b"0000000000000000_0000000000000000_0000011100110111_1100110000100000"; -- 0.028195150196552277
	pesos_i(3964) := b"1111111111111111_1111111111111111_1110111000000110_1000100111100000"; -- -0.07021272927522659
	pesos_i(3965) := b"0000000000000000_0000000000000000_0000100011111000_1110001011000000"; -- 0.03504769504070282
	pesos_i(3966) := b"0000000000000000_0000000000000000_0010010111100001_1110011011000000"; -- 0.14797823131084442
	pesos_i(3967) := b"1111111111111111_1111111111111111_1111111110010111_1011010000111101"; -- -0.0015914298128336668
	pesos_i(3968) := b"1111111111111111_1111111111111111_1111011101100001_0101110001010000"; -- -0.03367064520716667
	pesos_i(3969) := b"0000000000000000_0000000000000000_0000000101001000_1101001000000110"; -- 0.005017401184886694
	pesos_i(3970) := b"1111111111111111_1111111111111111_1111010110101001_1101110010100000"; -- -0.04037686437368393
	pesos_i(3971) := b"0000000000000000_0000000000000000_0001100101001010_0011100010000000"; -- 0.09878876805305481
	pesos_i(3972) := b"1111111111111111_1111111111111111_1101010011110101_1000101101000000"; -- -0.16812829673290253
	pesos_i(3973) := b"0000000000000000_0000000000000000_0101111100111111_1111001010000000"; -- 0.37206950783729553
	pesos_i(3974) := b"0000000000000000_0000000000000000_0011010110101010_0111111101000000"; -- 0.20963282883167267
	pesos_i(3975) := b"1111111111111111_1111111111111111_1101001101010100_0000101010000000"; -- -0.17449888586997986
	pesos_i(3976) := b"1111111111111111_1111111111111111_1101000011100101_0101111100000000"; -- -0.18400007486343384
	pesos_i(3977) := b"0000000000000000_0000000000000000_0010001101000000_0110011010000000"; -- 0.13770142197608948
	pesos_i(3978) := b"1111111111111111_1111111111111111_1010100110101011_1011111000000000"; -- -0.3372231721878052
	pesos_i(3979) := b"1111111111111111_1111111111111111_1100001010111010_1001100000000000"; -- -0.23934030532836914
	pesos_i(3980) := b"1111111111111111_1111111111111111_1111110101111100_0001101110100000"; -- -0.00982501357793808
	pesos_i(3981) := b"1111111111111111_1111111111111111_1111101000010100_0001000000000000"; -- -0.023131370544433594
	pesos_i(3982) := b"1111111111111111_1111111111111111_1101110101110100_0110010100000000"; -- -0.13494271039962769
	pesos_i(3983) := b"1111111111111111_1111111111111111_1110010111101001_1101001011000000"; -- -0.10190089046955109
	pesos_i(3984) := b"1111111111111111_1111111111111111_1111010001100001_1011110001010000"; -- -0.045383673161268234
	pesos_i(3985) := b"0000000000000000_0000000000000000_0010010101110111_0010111110000000"; -- 0.14634987711906433
	pesos_i(3986) := b"0000000000000000_0000000000000000_0011110100011111_0001001101000000"; -- 0.23875541985034943
	pesos_i(3987) := b"1111111111111111_1111111111111111_1110001110001100_1010000000100000"; -- -0.11113547533750534
	pesos_i(3988) := b"0000000000000000_0000000000000000_0010111001101101_0000000001000000"; -- 0.1813507229089737
	pesos_i(3989) := b"1111111111111111_1111111111111111_1100100111001010_1100100010000000"; -- -0.21174952387809753
	pesos_i(3990) := b"1111111111111111_1111111111111111_1111011110011011_0101001001000000"; -- -0.032786235213279724
	pesos_i(3991) := b"1111111111111111_1111111111111111_1111110111100101_0011011010001000"; -- -0.008221236988902092
	pesos_i(3992) := b"0000000000000000_0000000000000000_0001100011101110_1101100000000000"; -- 0.09739446640014648
	pesos_i(3993) := b"0000000000000000_0000000000000000_0000110011011110_1011011000000000"; -- 0.05027329921722412
	pesos_i(3994) := b"1111111111111111_1111111111111111_1111111010010000_0010111000011110"; -- -0.005612485576421022
	pesos_i(3995) := b"1111111111111111_1111111111111111_1011100100101000_0111010000000000"; -- -0.27672648429870605
	pesos_i(3996) := b"0000000000000000_0000000000000000_0011100000001000_1111100101000000"; -- 0.21888692677021027
	pesos_i(3997) := b"0000000000000000_0000000000000000_0010110000100111_0101010001000000"; -- 0.17247511446475983
	pesos_i(3998) := b"1111111111111111_1111111111111111_1011111011011010_1101011110000000"; -- -0.2544732391834259
	pesos_i(3999) := b"1111111111111111_1111111111111111_1111101011100001_0011111111110000"; -- -0.020000461488962173
	pesos_i(4000) := b"0000000000000000_0000000000000000_0011000001111000_1010000011000000"; -- 0.18934063613414764
	pesos_i(4001) := b"1111111111111111_1111111111111111_1010111110100101_0101011010000000"; -- -0.31388339400291443
	pesos_i(4002) := b"0000000000000000_0000000000000000_0001101001110110_1100011000100000"; -- 0.10337484627962112
	pesos_i(4003) := b"0000000000000000_0000000000000000_0010000100101110_0111011110000000"; -- 0.12961527705192566
	pesos_i(4004) := b"1111111111111111_1111111111111111_1111110101001001_0101011110011100"; -- -0.010599636472761631
	pesos_i(4005) := b"0000000000000000_0000000000000000_0001000011000111_1100011100100000"; -- 0.0655483677983284
	pesos_i(4006) := b"1111111111111111_1111111111111111_1111100111101011_1111100110101000"; -- -0.023743053898215294
	pesos_i(4007) := b"0000000000000000_0000000000000000_0001100101111000_0110011001100000"; -- 0.09949340671300888
	pesos_i(4008) := b"1111111111111111_1111111111111111_0111011100110010_1110011000000000"; -- -0.5343796014785767
	pesos_i(4009) := b"0000000000000000_0000000000000000_0010011000100010_0010011111000000"; -- 0.14895866811275482
	pesos_i(4010) := b"1111111111111111_1111111111111111_1110010000110010_0001001110000000"; -- -0.10861089825630188
	pesos_i(4011) := b"1111111111111111_1111111111111111_1001001110011011_0010111000000000"; -- -0.42341339588165283
	pesos_i(4012) := b"0000000000000000_0000000000000000_0010110101011011_1010111010000000"; -- 0.1771802008152008
	pesos_i(4013) := b"1111111111111111_1111111111111111_1101011111111111_0101001110000000"; -- -0.15626028180122375
	pesos_i(4014) := b"0000000000000000_0000000000000000_0011001111011001_0000100111000000"; -- 0.20253048837184906
	pesos_i(4015) := b"1111111111111111_1111111111111111_1110101010000100_1100111110000000"; -- -0.0839109718799591
	pesos_i(4016) := b"1111111111111111_1111111111111111_1111000010110100_0111000010010000"; -- -0.05974670872092247
	pesos_i(4017) := b"0000000000000000_0000000000000000_0000011001111111_1111101011011000"; -- 0.025390317663550377
	pesos_i(4018) := b"1111111111111111_1111111111111111_1100101011001001_0011001110000000"; -- -0.20786741375923157
	pesos_i(4019) := b"1111111111111111_1111111111111111_1111010101110111_1000110011000000"; -- -0.041144564747810364
	pesos_i(4020) := b"0000000000000000_0000000000000000_0010111010101011_0100001001000000"; -- 0.18230070173740387
	pesos_i(4021) := b"0000000000000000_0000000000000000_0000110110001100_1011100011000000"; -- 0.05292849242687225
	pesos_i(4022) := b"0000000000000000_0000000000000000_0011010100000110_0110000111000000"; -- 0.2071286290884018
	pesos_i(4023) := b"1111111111111111_1111111111111111_1101100001001000_0110101000000000"; -- -0.1551450490951538
	pesos_i(4024) := b"1111111111111111_1111111111111111_1110001110010010_1111100001100000"; -- -0.11103866249322891
	pesos_i(4025) := b"1111111111111111_1111111111111111_1100101111011110_1110110100000000"; -- -0.20362967252731323
	pesos_i(4026) := b"1111111111111111_1111111111111111_1011101111111000_1001111100000000"; -- -0.2657375931739807
	pesos_i(4027) := b"1111111111111111_1111111111111111_1110010011000111_0100010111000000"; -- -0.10633434355258942
	pesos_i(4028) := b"0000000000000000_0000000000000000_0001010000100111_1110010011100000"; -- 0.07873373478651047
	pesos_i(4029) := b"0000000000000000_0000000000000000_0001100111101010_1101110011100000"; -- 0.10123997181653976
	pesos_i(4030) := b"1111111111111111_1111111111111111_1011001011011000_1010000100000000"; -- -0.30138200521469116
	pesos_i(4031) := b"0000000000000000_0000000000000000_0010001011101000_0001011110000000"; -- 0.13635393977165222
	pesos_i(4032) := b"1111111111111111_1111111111111111_1001000101101101_1001110100000000"; -- -0.43192118406295776
	pesos_i(4033) := b"0000000000000000_0000000000000000_0011010101001001_1100110110000000"; -- 0.20815739035606384
	pesos_i(4034) := b"0000000000000000_0000000000000000_0010010101101100_1011101011000000"; -- 0.1461903303861618
	pesos_i(4035) := b"1111111111111111_1111111111111111_1110110111011100_1101000110100000"; -- -0.07084932178258896
	pesos_i(4036) := b"1111111111111111_1111111111111111_1100101011111101_0011001110000000"; -- -0.20707395672798157
	pesos_i(4037) := b"1111111111111111_1111111111111111_1111100011111010_0100110110111000"; -- -0.027430670335888863
	pesos_i(4038) := b"0000000000000000_0000000000000000_0011000010110000_1101001000000000"; -- 0.19019806385040283
	pesos_i(4039) := b"0000000000000000_0000000000000000_0000001001011010_1010010101001100"; -- 0.009195643477141857
	pesos_i(4040) := b"1111111111111111_1111111111111111_1101000101010000_0101010010000000"; -- -0.18236801028251648
	pesos_i(4041) := b"1111111111111111_1111111111111111_1101011111110010_0111010000000000"; -- -0.15645670890808105
	pesos_i(4042) := b"1111111111111111_1111111111111111_1101001100110110_1011010111000000"; -- -0.17494644224643707
	pesos_i(4043) := b"1111111111111111_1111111111111111_1110010101000100_1000010110100000"; -- -0.10442318767309189
	pesos_i(4044) := b"0000000000000000_0000000000000000_0011011101101001_0111011100000000"; -- 0.21645301580429077
	pesos_i(4045) := b"1111111111111111_1111111111111111_1111101001101010_0000101101101000"; -- -0.02181938849389553
	pesos_i(4046) := b"1111111111111111_1111111111111111_1101010101110010_1110011010000000"; -- -0.16621550917625427
	pesos_i(4047) := b"1111111111111111_1111111111111111_1100010011000110_1000011010000000"; -- -0.2313457429409027
	pesos_i(4048) := b"1111111111111111_1111111111111111_1101000011000110_0101001001000000"; -- -0.18447385728359222
	pesos_i(4049) := b"1111111111111111_1111111111111111_0101111100101111_0000101100000000"; -- -0.62818843126297
	pesos_i(4050) := b"0000000000000000_0000000000000000_0000110010001111_1011110111000000"; -- 0.04906831681728363
	pesos_i(4051) := b"0000000000000000_0000000000000000_0001111001110011_0011101010000000"; -- 0.11894574761390686
	pesos_i(4052) := b"0000000000000000_0000000000000000_0001110011011101_1000001110100000"; -- 0.11275503784418106
	pesos_i(4053) := b"1111111111111111_1111111111111111_1111001100111110_0001100100000000"; -- -0.049833714962005615
	pesos_i(4054) := b"0000000000000000_0000000000000000_0000010100010110_1100001001000000"; -- 0.01987852156162262
	pesos_i(4055) := b"1111111111111111_1111111111111111_1101111101010001_1010110101000000"; -- -0.12765996158123016
	pesos_i(4056) := b"0000000000000000_0000000000000000_0000001000010110_0001100011011100"; -- 0.008149675093591213
	pesos_i(4057) := b"1111111111111111_1111111111111111_1110010110001110_0011101101000000"; -- -0.10329847037792206
	pesos_i(4058) := b"1111111111111111_1111111111111111_0110000001001101_1000101000000000"; -- -0.6238168478012085
	pesos_i(4059) := b"1111111111111111_1111111111111111_1101010010111111_1000101100000000"; -- -0.16895228624343872
	pesos_i(4060) := b"0000000000000000_0000000000000000_0000000011001000_1000111001010010"; -- 0.003060240764170885
	pesos_i(4061) := b"1111111111111111_1111111111111111_1100011001110111_1111100000000000"; -- -0.2247319221496582
	pesos_i(4062) := b"1111111111111111_1111111111111111_1110100010001101_0000001010100000"; -- -0.09159835427999496
	pesos_i(4063) := b"1111111111111111_1111111111111111_1101001100110111_0101100001000000"; -- -0.17493675649166107
	pesos_i(4064) := b"0000000000000000_0000000000000000_0010110011010000_0001101001000000"; -- 0.17505039274692535
	pesos_i(4065) := b"0000000000000000_0000000000000000_0000100111111110_1111100101010000"; -- 0.039046842604875565
	pesos_i(4066) := b"1111111111111111_1111111111111111_1111101110101000_1001000001000000"; -- -0.01695917546749115
	pesos_i(4067) := b"1111111111111111_1111111111111111_1010111001100001_1100010110000000"; -- -0.31882062554359436
	pesos_i(4068) := b"1111111111111111_1111111111111111_1101110011000011_1011000110000000"; -- -0.13763895630836487
	pesos_i(4069) := b"0000000000000000_0000000000000000_0010011100010111_0100001010000000"; -- 0.15269866585731506
	pesos_i(4070) := b"0000000000000000_0000000000000000_0100100000011111_1111111100000000"; -- 0.2817382216453552
	pesos_i(4071) := b"1111111111111111_1111111111111111_1001111110111111_1100110000000000"; -- -0.3759796619415283
	pesos_i(4072) := b"1111111111111111_1111111111111111_1101111111110110_0000001011000000"; -- -0.12515242397785187
	pesos_i(4073) := b"1111111111111111_1111111111111111_1000011011101101_0000011110000000"; -- -0.4729457199573517
	pesos_i(4074) := b"1111111111111111_1111111111111111_1010110111101110_0001000010000000"; -- -0.3205861747264862
	pesos_i(4075) := b"0000000000000000_0000000000000000_0100101111001100_1001101110000000"; -- 0.2960908114910126
	pesos_i(4076) := b"1111111111111111_1111111111111111_1010000101010111_1011100110000000"; -- -0.36975517868995667
	pesos_i(4077) := b"1111111111111111_1111111111111111_1111100111000100_0100101101100000"; -- -0.024348534643650055
	pesos_i(4078) := b"1111111111111111_1111111111111111_1110110110011100_0010000010100000"; -- -0.0718364343047142
	pesos_i(4079) := b"1111111111111111_1111111111111111_1101000001100011_1010010100000000"; -- -0.18597954511642456
	pesos_i(4080) := b"0000000000000000_0000000000000000_0011000010101111_0111001011000000"; -- 0.19017712771892548
	pesos_i(4081) := b"0000000000000000_0000000000000000_0110100000110101_1100111110000000"; -- 0.4070710837841034
	pesos_i(4082) := b"1111111111111111_1111111111111111_1110011110100110_0011100010000000"; -- -0.09511992335319519
	pesos_i(4083) := b"1111111111111111_1111111111111111_1011000111011101_0101000110000000"; -- -0.3052166998386383
	pesos_i(4084) := b"1111111111111111_1111111111111111_1111111111101101_0010010100000111"; -- -0.00028770993230864406
	pesos_i(4085) := b"1111111111111111_1111111111111111_1010111100011101_1000111010000000"; -- -0.315955251455307
	pesos_i(4086) := b"1111111111111111_1111111111111111_1010000101000101_0111101010000000"; -- -0.3700335919857025
	pesos_i(4087) := b"1111111111111111_1111111111111111_1000110110110010_0101101100000000"; -- -0.44649726152420044
	pesos_i(4088) := b"1111111111111111_1111111111111111_1011110000001110_0111011000000000"; -- -0.2654043436050415
	pesos_i(4089) := b"1111111111111111_1111111111111111_1111110001011010_1111101101101000"; -- -0.014236724004149437
	pesos_i(4090) := b"1111111111111111_1111111111111111_1101111101101011_1001011110000000"; -- -0.12726452946662903
	pesos_i(4091) := b"1111111111111111_1111111111111111_1100000101010011_0100110110000000"; -- -0.2448226511478424
	pesos_i(4092) := b"0000000000000000_0000000000000000_0010100001111101_0001101000000000"; -- 0.15815889835357666
	pesos_i(4093) := b"1111111111111111_1111111111111111_0101010001100011_1101001100000000"; -- -0.6703518033027649
	pesos_i(4094) := b"0000000000000000_0000000000000000_0001100110011100_0110001011100000"; -- 0.10004251450300217
	pesos_i(4095) := b"1111111111111111_1111111111111111_1011100111000010_1000001100000000"; -- -0.2743757367134094
	pesos_i(4096) := b"0000000000000000_0000000000000000_0001111000101010_0101001000100000"; -- 0.11783326417207718
	pesos_i(4097) := b"0000000000000000_0000000000000000_0110011011101010_0100110000000000"; -- 0.40201258659362793
	pesos_i(4098) := b"1111111111111111_1111111111111111_1011110001001101_1001010010000000"; -- -0.26444122195243835
	pesos_i(4099) := b"1111111111111111_1111111111111111_1100000010010010_1111011010000000"; -- -0.24775752425193787
	pesos_i(4100) := b"0000000000000000_0000000000000000_0101010100101110_0000100010000000"; -- 0.3327336609363556
	pesos_i(4101) := b"1111111111111111_1111111111111111_1111001111011100_0100011100110000"; -- -0.04742007330060005
	pesos_i(4102) := b"0000000000000000_0000000000000000_0001001100001101_0001100011000000"; -- 0.07441858947277069
	pesos_i(4103) := b"1111111111111111_1111111111111111_1110001011101000_0101101011000000"; -- -0.11364205181598663
	pesos_i(4104) := b"0000000000000000_0000000000000000_0001110011100000_0111011110000000"; -- 0.11280009150505066
	pesos_i(4105) := b"1111111111111111_1111111111111111_1101110010110001_1111011101000000"; -- -0.13790945708751678
	pesos_i(4106) := b"0000000000000000_0000000000000000_0100110101001010_1011000000000000"; -- 0.30192089080810547
	pesos_i(4107) := b"0000000000000000_0000000000000000_0001000101010100_1000101100100000"; -- 0.06769628077745438
	pesos_i(4108) := b"1111111111111111_1111111111111111_1101010100000101_0111000001000000"; -- -0.16788576543331146
	pesos_i(4109) := b"1111111111111111_1111111111111111_1100110110100011_1100010111000000"; -- -0.19671978056430817
	pesos_i(4110) := b"1111111111111111_1111111111111111_1101000111111101_1111100011000000"; -- -0.17971844971179962
	pesos_i(4111) := b"1111111111111111_1111111111111111_1110110010100010_1111100110000000"; -- -0.07563820481300354
	pesos_i(4112) := b"0000000000000000_0000000000000000_0001001010100100_0010010011000000"; -- 0.0728171318769455
	pesos_i(4113) := b"1111111111111111_1111111111111111_1111010001001010_1101010001110000"; -- -0.04573318734765053
	pesos_i(4114) := b"1111111111111111_1111111111111111_1110111100010010_1111101011000000"; -- -0.06611664593219757
	pesos_i(4115) := b"1111111111111111_1111111111111111_1011000111010111_1000001100000000"; -- -0.3053053021430969
	pesos_i(4116) := b"1111111111111111_1111111111111111_1110000100110010_0101111111100000"; -- -0.12032509595155716
	pesos_i(4117) := b"0000000000000000_0000000000000000_0011011001011011_0001011010000000"; -- 0.21232739090919495
	pesos_i(4118) := b"1111111111111111_1111111111111111_1110011010110100_1011001000100000"; -- -0.09880530089139938
	pesos_i(4119) := b"1111111111111111_1111111111111111_1110101101010011_0101100110000000"; -- -0.0807594358921051
	pesos_i(4120) := b"0000000000000000_0000000000000000_0001010001110111_1100111110100000"; -- 0.07995317131280899
	pesos_i(4121) := b"1111111111111111_1111111111111111_1101011100000010_1111110001000000"; -- -0.1601106971502304
	pesos_i(4122) := b"0000000000000000_0000000000000000_0010111010111011_1001110010000000"; -- 0.18255022168159485
	pesos_i(4123) := b"1111111111111111_1111111111111111_1011110110010111_1000100010000000"; -- -0.25940653681755066
	pesos_i(4124) := b"0000000000000000_0000000000000000_0000111100111010_0101000000100000"; -- 0.05948353558778763
	pesos_i(4125) := b"1111111111111111_1111111111111111_1010100110010001_1010011110000000"; -- -0.3376212418079376
	pesos_i(4126) := b"0000000000000000_0000000000000000_0011110011111000_1000011110000000"; -- 0.23816725611686707
	pesos_i(4127) := b"1111111111111111_1111111111111111_1110110000101010_0100001001100000"; -- -0.07748017460107803
	pesos_i(4128) := b"0000000000000000_0000000000000000_0011010100101001_0010111001000000"; -- 0.20765961706638336
	pesos_i(4129) := b"0000000000000000_0000000000000000_0001001111111000_0011101110100000"; -- 0.07800648361444473
	pesos_i(4130) := b"0000000000000000_0000000000000000_0001000101001011_1000110011100000"; -- 0.06755905598402023
	pesos_i(4131) := b"1111111111111111_1111111111111111_1110110110000101_0000111000000000"; -- -0.07218849658966064
	pesos_i(4132) := b"0000000000000000_0000000000000000_0001110110011010_0001100110100000"; -- 0.11563263088464737
	pesos_i(4133) := b"0000000000000000_0000000000000000_0001110100001110_1111011111000000"; -- 0.1135096400976181
	pesos_i(4134) := b"1111111111111111_1111111111111111_1110110001111100_1010100010000000"; -- -0.07622286677360535
	pesos_i(4135) := b"1111111111111111_1111111111111111_1111111010000100_0111001001001010"; -- -0.005791527684777975
	pesos_i(4136) := b"1111111111111111_1111111111111111_1100111110111001_0100101000000000"; -- -0.18857896327972412
	pesos_i(4137) := b"0000000000000000_0000000000000000_0001000110111001_1000011111100000"; -- 0.06923722475767136
	pesos_i(4138) := b"1111111111111111_1111111111111111_1101000011110110_0001101111000000"; -- -0.18374468386173248
	pesos_i(4139) := b"1111111111111111_1111111111111111_1110011010111101_0111101001000000"; -- -0.09867130219936371
	pesos_i(4140) := b"1111111111111111_1111111111111111_1101111110101011_1100110100000000"; -- -0.12628477811813354
	pesos_i(4141) := b"1111111111111111_1111111111111111_1100110100110001_0101100110000000"; -- -0.1984657347202301
	pesos_i(4142) := b"0000000000000000_0000000000000000_0011000011001011_1101011000000000"; -- 0.19061028957366943
	pesos_i(4143) := b"1111111111111111_1111111111111111_1111010110100111_1000101011100000"; -- -0.04041225463151932
	pesos_i(4144) := b"0000000000000000_0000000000000000_0010011010111001_1110001011000000"; -- 0.15127389132976532
	pesos_i(4145) := b"1111111111111111_1111111111111111_1011011010011010_0001111110000000"; -- -0.2867107689380646
	pesos_i(4146) := b"1111111111111111_1111111111111111_1100110001010011_1001111101000000"; -- -0.20184902846813202
	pesos_i(4147) := b"0000000000000000_0000000000000000_0100011111111111_1001111110000000"; -- 0.2812442481517792
	pesos_i(4148) := b"1111111111111111_1111111111111111_1110101001101011_1010001000100000"; -- -0.08429514616727829
	pesos_i(4149) := b"0000000000000000_0000000000000000_0001001101101110_1110111011100000"; -- 0.07591145485639572
	pesos_i(4150) := b"0000000000000000_0000000000000000_0001000101100111_0001010111100000"; -- 0.06797920912504196
	pesos_i(4151) := b"0000000000000000_0000000000000000_0010111011101110_0111000010000000"; -- 0.18332579731941223
	pesos_i(4152) := b"0000000000000000_0000000000000000_0010000101001010_0001001111000000"; -- 0.13003657758235931
	pesos_i(4153) := b"1111111111111111_1111111111111111_1111100110000110_0001010001010000"; -- -0.025297861546278
	pesos_i(4154) := b"0000000000000000_0000000000000000_0000111010001101_1100001101110000"; -- 0.05685063824057579
	pesos_i(4155) := b"0000000000000000_0000000000000000_0001111100111101_0001000001000000"; -- 0.1220255047082901
	pesos_i(4156) := b"0000000000000000_0000000000000000_0010011011100101_0001100001000000"; -- 0.1519332081079483
	pesos_i(4157) := b"1111111111111111_1111111111111111_1011110111000101_0010000110000000"; -- -0.2587107717990875
	pesos_i(4158) := b"0000000000000000_0000000000000000_0000011100111001_1001100011100000"; -- 0.028222613036632538
	pesos_i(4159) := b"1111111111111111_1111111111111111_1100000000100011_1100011010000000"; -- -0.24945411086082458
	pesos_i(4160) := b"0000000000000000_0000000000000000_0011000110010011_1111110110000000"; -- 0.19366440176963806
	pesos_i(4161) := b"0000000000000000_0000000000000000_0011111011010001_0000001110000000"; -- 0.2453767955303192
	pesos_i(4162) := b"1111111111111111_1111111111111111_1111111011111110_0110011011010100"; -- -0.0039306385442614555
	pesos_i(4163) := b"0000000000000000_0000000000000000_0001001010001111_1111010111100000"; -- 0.07250916212797165
	pesos_i(4164) := b"0000000000000000_0000000000000000_0010001111000000_0001000011000000"; -- 0.1396494358778
	pesos_i(4165) := b"1111111111111111_1111111111111111_1100110010000011_1100101111000000"; -- -0.20111395418643951
	pesos_i(4166) := b"1111111111111111_1111111111111111_1101110010100111_0100110111000000"; -- -0.1380721479654312
	pesos_i(4167) := b"0000000000000000_0000000000000000_0001000010000010_0111110001100000"; -- 0.06449105590581894
	pesos_i(4168) := b"0000000000000000_0000000000000000_0011100000101001_1110010000000000"; -- 0.2193892002105713
	pesos_i(4169) := b"1111111111111111_1111111111111111_1101101111111110_0011000001000000"; -- -0.1406526416540146
	pesos_i(4170) := b"1111111111111111_1111111111111111_1111110101001010_1100111100001100"; -- -0.01057725865393877
	pesos_i(4171) := b"0000000000000000_0000000000000000_0001001001111000_0000010000100000"; -- 0.0721438005566597
	pesos_i(4172) := b"1111111111111111_1111111111111111_1110110111001111_0001010111000000"; -- -0.07105888426303864
	pesos_i(4173) := b"0000000000000000_0000000000000000_0001000001010010_1100011100000000"; -- 0.0637630820274353
	pesos_i(4174) := b"1111111111111111_1111111111111111_1010111100001100_1101000110000000"; -- -0.31621065735816956
	pesos_i(4175) := b"0000000000000000_0000000000000000_0010011011001000_1010010011000000"; -- 0.15149907767772675
	pesos_i(4176) := b"1111111111111111_1111111111111111_1111011111000111_0000010000010000"; -- -0.0321195088326931
	pesos_i(4177) := b"0000000000000000_0000000000000000_0101011001111111_0110011110000000"; -- 0.33788153529167175
	pesos_i(4178) := b"1111111111111111_1111111111111111_1110001000101011_0000110110100000"; -- -0.11653055995702744
	pesos_i(4179) := b"1111111111111111_1111111111111111_1100101111000000_0100111011000000"; -- -0.20409686863422394
	pesos_i(4180) := b"0000000000000000_0000000000000000_0000001010000011_1100111010000100"; -- 0.009823710657656193
	pesos_i(4181) := b"0000000000000000_0000000000000000_0001101111000101_1111111110100000"; -- 0.10848996788263321
	pesos_i(4182) := b"1111111111111111_1111111111111111_1111011011111010_1001101110010000"; -- -0.03523853048682213
	pesos_i(4183) := b"1111111111111111_1111111111111111_1100000100010100_0011110010000000"; -- -0.2457849681377411
	pesos_i(4184) := b"0000000000000000_0000000000000000_0010100100010100_0110100010000000"; -- 0.16046765446662903
	pesos_i(4185) := b"1111111111111111_1111111111111111_1101111100000100_0110111001000000"; -- -0.1288386434316635
	pesos_i(4186) := b"1111111111111111_1111111111111111_1111100111110011_0101110011010000"; -- -0.023630332201719284
	pesos_i(4187) := b"1111111111111111_1111111111111111_1101011010111010_0000101011000000"; -- -0.16122372448444366
	pesos_i(4188) := b"1111111111111111_1111111111111111_1101111011110111_1110011000000000"; -- -0.12902987003326416
	pesos_i(4189) := b"1111111111111111_1111111111111111_1111011011111011_0110011000000000"; -- -0.03522646427154541
	pesos_i(4190) := b"1111111111111111_1111111111111111_1101011000110110_1010111111000000"; -- -0.16322804987430573
	pesos_i(4191) := b"0000000000000000_0000000000000000_0000100000010110_1100100000100000"; -- 0.031597621738910675
	pesos_i(4192) := b"0000000000000000_0000000000000000_0010111100010000_0110001100000000"; -- 0.18384379148483276
	pesos_i(4193) := b"0000000000000000_0000000000000000_0010000001000111_0101101010000000"; -- 0.12608876824378967
	pesos_i(4194) := b"0000000000000000_0000000000000000_0000101011011010_1111010011010000"; -- 0.042403507977724075
	pesos_i(4195) := b"1111111111111111_1111111111111111_1101101101010111_1000110100000000"; -- -0.14319533109664917
	pesos_i(4196) := b"0000000000000000_0000000000000000_0001011010010001_1001000110100000"; -- 0.08815870434045792
	pesos_i(4197) := b"0000000000000000_0000000000000000_0001111111111001_1101100110000000"; -- 0.12490615248680115
	pesos_i(4198) := b"1111111111111111_1111111111111111_1111110010001010_0001101100010000"; -- -0.013517674058675766
	pesos_i(4199) := b"0000000000000000_0000000000000000_0000100000001000_1100111100110000"; -- 0.0313844196498394
	pesos_i(4200) := b"1111111111111111_1111111111111111_1111001001100000_1000100111110000"; -- -0.053214434534311295
	pesos_i(4201) := b"0000000000000000_0000000000000000_0000101100011010_0011111011100000"; -- 0.04336922615766525
	pesos_i(4202) := b"1111111111111111_1111111111111111_1111001111001001_0010110111100000"; -- -0.04771149903535843
	pesos_i(4203) := b"0000000000000000_0000000000000000_0001000000110011_1101111000000000"; -- 0.06329143047332764
	pesos_i(4204) := b"0000000000000000_0000000000000000_0011110110101100_1111101011000000"; -- 0.24092070758342743
	pesos_i(4205) := b"1111111111111111_1111111111111111_1011110101010110_0001011110000000"; -- -0.2604050934314728
	pesos_i(4206) := b"1111111111111111_1111111111111111_1011100010100111_1100010010000000"; -- -0.27869006991386414
	pesos_i(4207) := b"1111111111111111_1111111111111111_1010111010100011_1100100000000000"; -- -0.3178133964538574
	pesos_i(4208) := b"0000000000000000_0000000000000000_0001000101010010_1000001101000000"; -- 0.06766529381275177
	pesos_i(4209) := b"0000000000000000_0000000000000000_0010000101110001_0010101001000000"; -- 0.13063301146030426
	pesos_i(4210) := b"0000000000000000_0000000000000000_0000100010011110_1110001100010000"; -- 0.03367442265152931
	pesos_i(4211) := b"0000000000000000_0000000000000000_0001111100100011_1011011110000000"; -- 0.12163874506950378
	pesos_i(4212) := b"1111111111111111_1111111111111111_1101101010101011_0101111010000000"; -- -0.14582261443138123
	pesos_i(4213) := b"1111111111111111_1111111111111111_1101100110100111_0101100111000000"; -- -0.1497901827096939
	pesos_i(4214) := b"0000000000000000_0000000000000000_0000110010110100_0111110100110000"; -- 0.04962904378771782
	pesos_i(4215) := b"0000000000000000_0000000000000000_0010000001101011_1000010000000000"; -- 0.12664055824279785
	pesos_i(4216) := b"1111111111111111_1111111111111111_1110111100110010_1111001001100000"; -- -0.06562886387109756
	pesos_i(4217) := b"0000000000000000_0000000000000000_0000110000101010_1010010001000000"; -- 0.04752565920352936
	pesos_i(4218) := b"1111111111111111_1111111111111111_1110111001111000_1111111000100000"; -- -0.06846629828214645
	pesos_i(4219) := b"0000000000000000_0000000000000000_0001111111000101_1110111001100000"; -- 0.12411393970251083
	pesos_i(4220) := b"1111111111111111_1111111111111111_1110111001000011_0100000110000000"; -- -0.06928625702857971
	pesos_i(4221) := b"1111111111111111_1111111111111111_1110001100111001_0100011000000000"; -- -0.11240732669830322
	pesos_i(4222) := b"1111111111111111_1111111111111111_1111011001110100_0010010011100000"; -- -0.03729028254747391
	pesos_i(4223) := b"0000000000000000_0000000000000000_0100000111010010_0010001100000000"; -- 0.25711268186569214
	pesos_i(4224) := b"1111111111111111_1111111111111111_1110010101011101_0010000010000000"; -- -0.1040477454662323
	pesos_i(4225) := b"1111111111111111_1111111111111111_1100010001100000_1001001010000000"; -- -0.2329014241695404
	pesos_i(4226) := b"1111111111111111_1111111111111111_1110001011010111_1010110011100000"; -- -0.11389655619859695
	pesos_i(4227) := b"0000000000000000_0000000000000000_0000010110010110_1001111000111000"; -- 0.021829498931765556
	pesos_i(4228) := b"1111111111111111_1111111111111111_1110110011011000_1010010100000000"; -- -0.07481926679611206
	pesos_i(4229) := b"0000000000000000_0000000000000000_0011110110001011_0100010001000000"; -- 0.24040628969669342
	pesos_i(4230) := b"1111111111111111_1111111111111111_1110101100111010_0011111011100000"; -- -0.08114249259233475
	pesos_i(4231) := b"0000000000000000_0000000000000000_0010100001111000_0111001110000000"; -- 0.15808793902397156
	pesos_i(4232) := b"0000000000000000_0000000000000000_0001110000101101_0110111010000000"; -- 0.11006823182106018
	pesos_i(4233) := b"0000000000000000_0000000000000000_0000010001000101_1111000111001000"; -- 0.0166922677308321
	pesos_i(4234) := b"0000000000000000_0000000000000000_0100000000010010_0110011010000000"; -- 0.2502807676792145
	pesos_i(4235) := b"1111111111111111_1111111111111111_1111111111110110_1100101101100100"; -- -0.00014046498108655214
	pesos_i(4236) := b"0000000000000000_0000000000000000_0001100001101010_0000011000100000"; -- 0.09536779671907425
	pesos_i(4237) := b"1111111111111111_1111111111111111_1101110000001101_1100010111000000"; -- -0.14041484892368317
	pesos_i(4238) := b"0000000000000000_0000000000000000_0001111001111001_0000100101100000"; -- 0.11903437227010727
	pesos_i(4239) := b"0000000000000000_0000000000000000_0000110000010010_0101000001000000"; -- 0.047154441475868225
	pesos_i(4240) := b"0000000000000000_0000000000000000_0100011100111011_0111111100000000"; -- 0.278251588344574
	pesos_i(4241) := b"1111111111111111_1111111111111111_1110001001000100_1100001101000000"; -- -0.1161382645368576
	pesos_i(4242) := b"0000000000000000_0000000000000000_0000111010100100_1011010100000000"; -- 0.057200729846954346
	pesos_i(4243) := b"0000000000000000_0000000000000000_0000110000101110_0101101110010000"; -- 0.04758236184716225
	pesos_i(4244) := b"1111111111111111_1111111111111111_1101100001110111_0011001001000000"; -- -0.15443120896816254
	pesos_i(4245) := b"0000000000000000_0000000000000000_0011110001111100_0010000101000000"; -- 0.23626907169818878
	pesos_i(4246) := b"1111111111111111_1111111111111111_1110111100001001_1110110011000000"; -- -0.06625480949878693
	pesos_i(4247) := b"0000000000000000_0000000000000000_0010000110000110_1000000011000000"; -- 0.13095860183238983
	pesos_i(4248) := b"0000000000000000_0000000000000000_0100010101111110_0011000110000000"; -- 0.2714568078517914
	pesos_i(4249) := b"0000000000000000_0000000000000000_0001110010101101_1001110100100000"; -- 0.11202413588762283
	pesos_i(4250) := b"0000000000000000_0000000000000000_0010001010000001_1100101001000000"; -- 0.13479293882846832
	pesos_i(4251) := b"1111111111111111_1111111111111111_1101010000110001_1101110101000000"; -- -0.17111413180828094
	pesos_i(4252) := b"0000000000000000_0000000000000000_0010101101010010_1111100101000000"; -- 0.16923482716083527
	pesos_i(4253) := b"1111111111111111_1111111111111111_1111101001011110_1101001011110000"; -- -0.02199060097336769
	pesos_i(4254) := b"1111111111111111_1111111111111111_1011110001110001_1100100010000000"; -- -0.26388880610466003
	pesos_i(4255) := b"0000000000000000_0000000000000000_0001110111010001_1100001000000000"; -- 0.11648190021514893
	pesos_i(4256) := b"0000000000000000_0000000000000000_0011001011011010_1100001001000000"; -- 0.19865049421787262
	pesos_i(4257) := b"0000000000000000_0000000000000000_0100111101001110_1111100110000000"; -- 0.30979880690574646
	pesos_i(4258) := b"0000000000000000_0000000000000000_0001101001110011_0100000101000000"; -- 0.1033211499452591
	pesos_i(4259) := b"1111111111111111_1111111111111111_1101100101011110_1100110000000000"; -- -0.15089726448059082
	pesos_i(4260) := b"1111111111111111_1111111111111111_1101001110011010_1100100001000000"; -- -0.17341946065425873
	pesos_i(4261) := b"1111111111111111_1111111111111111_1101100001000101_1010011111000000"; -- -0.15518714487552643
	pesos_i(4262) := b"1111111111111111_1111111111111111_1001011101110101_1000111010000000"; -- -0.408362478017807
	pesos_i(4263) := b"0000000000000000_0000000000000000_0100000000000000_1110010110000000"; -- 0.25001367926597595
	pesos_i(4264) := b"1111111111111111_1111111111111111_1101101100101100_0000000100000000"; -- -0.14385980367660522
	pesos_i(4265) := b"0000000000000000_0000000000000000_0001100000001100_0011001001000000"; -- 0.09393610060214996
	pesos_i(4266) := b"1111111111111111_1111111111111111_1110000011100001_0100111010100000"; -- -0.12156208604574203
	pesos_i(4267) := b"1111111111111111_1111111111111111_1101100001000111_1011101110000000"; -- -0.15515545010566711
	pesos_i(4268) := b"1111111111111111_1111111111111111_1100100011011100_0001001100000000"; -- -0.21539193391799927
	pesos_i(4269) := b"1111111111111111_1111111111111111_1111011110011001_0101010011000000"; -- -0.032816603779792786
	pesos_i(4270) := b"0000000000000000_0000000000000000_0010000111000010_1101110010000000"; -- 0.13187959790229797
	pesos_i(4271) := b"1111111111111111_1111111111111111_1010011000101000_1001100100000000"; -- -0.35094302892684937
	pesos_i(4272) := b"1111111111111111_1111111111111111_1110000110010011_1010010000000000"; -- -0.11884093284606934
	pesos_i(4273) := b"1111111111111111_1111111111111111_1011110110011000_0001101110000000"; -- -0.2593977749347687
	pesos_i(4274) := b"1111111111111111_1111111111111111_1001110011000001_1000001010000000"; -- -0.3876722753047943
	pesos_i(4275) := b"1111111111111111_1111111111111111_1110110111111111_1100111000000000"; -- -0.07031548023223877
	pesos_i(4276) := b"0000000000000000_0000000000000000_0011010011101110_1000101001000000"; -- 0.2067648321390152
	pesos_i(4277) := b"1111111111111111_1111111111111111_1100001001011111_0011000011000000"; -- -0.2407350093126297
	pesos_i(4278) := b"1111111111111111_1111111111111111_1001111111100001_1011011010000000"; -- -0.375462144613266
	pesos_i(4279) := b"0000000000000000_0000000000000000_0000000111101001_1010001101000100"; -- 0.007471279241144657
	pesos_i(4280) := b"0000000000000000_0000000000000000_0000110000000010_1011110101010000"; -- 0.04691680148243904
	pesos_i(4281) := b"1111111111111111_1111111111111111_1001000010000111_0010100110000000"; -- -0.4354375898838043
	pesos_i(4282) := b"1111111111111111_1111111111111111_1111100101001001_0001010000000000"; -- -0.026228666305541992
	pesos_i(4283) := b"1111111111111111_1111111111111111_1111101000101000_0011001110100000"; -- -0.02282407134771347
	pesos_i(4284) := b"0000000000000000_0000000000000000_0001100010111100_1010100110000000"; -- 0.09662875533103943
	pesos_i(4285) := b"1111111111111111_1111111111111111_1111101011111011_0010011100100000"; -- -0.019605211913585663
	pesos_i(4286) := b"0000000000000000_0000000000000000_0000001010111110_0000101100111000"; -- 0.010712338611483574
	pesos_i(4287) := b"1111111111111111_1111111111111111_1101100011000011_0110101110000000"; -- -0.15326812863349915
	pesos_i(4288) := b"0000000000000000_0000000000000000_0010011000100011_1101001011000000"; -- 0.1489841192960739
	pesos_i(4289) := b"1111111111111111_1111111111111111_1111111001011010_0111011011001110"; -- -0.006432127673178911
	pesos_i(4290) := b"1111111111111111_1111111111111111_1111110000101001_1001101100011100"; -- -0.014990144409239292
	pesos_i(4291) := b"0000000000000000_0000000000000000_0010001100100010_1111001010000000"; -- 0.13725200295448303
	pesos_i(4292) := b"0000000000000000_0000000000000000_0100001000110101_0110110110000000"; -- 0.2586277425289154
	pesos_i(4293) := b"1111111111111111_1111111111111111_1101110111101110_0001111010000000"; -- -0.13308534026145935
	pesos_i(4294) := b"1111111111111111_1111111111111111_1111011000101010_0111111110100000"; -- -0.03841402381658554
	pesos_i(4295) := b"1111111111111111_1111111111111111_1101011111100001_0110111101000000"; -- -0.15671639144420624
	pesos_i(4296) := b"0000000000000000_0000000000000000_0100000000001001_0100010100000000"; -- 0.250141441822052
	pesos_i(4297) := b"1111111111111111_1111111111111111_1110011010011001_0111100111000000"; -- -0.0992206484079361
	pesos_i(4298) := b"1111111111111111_1111111111111111_1101011111101011_0011111101000000"; -- -0.15656666457653046
	pesos_i(4299) := b"0000000000000000_0000000000000000_0001000100000001_1110100110000000"; -- 0.06643542647361755
	pesos_i(4300) := b"1111111111111111_1111111111111111_1100111110001101_0000101111000000"; -- -0.1892540603876114
	pesos_i(4301) := b"0000000000000000_0000000000000000_0001101001000001_1110001100000000"; -- 0.10256785154342651
	pesos_i(4302) := b"1111111111111111_1111111111111111_1101101011000010_1111011000000000"; -- -0.14546263217926025
	pesos_i(4303) := b"1111111111111111_1111111111111111_1011100011111101_1101000110000000"; -- -0.27737703919410706
	pesos_i(4304) := b"0000000000000000_0000000000000000_0001001010011011_1111000001100000"; -- 0.07269193977117538
	pesos_i(4305) := b"1111111111111111_1111111111111111_1100000111010010_0001101010000000"; -- -0.24288782477378845
	pesos_i(4306) := b"0000000000000000_0000000000000000_0000010111011000_0000001101000000"; -- 0.02282734215259552
	pesos_i(4307) := b"1111111111111111_1111111111111111_1111010100000100_0011000010110000"; -- -0.0429048128426075
	pesos_i(4308) := b"1111111111111111_1111111111111111_1010110110101011_1100010100000000"; -- -0.32159775495529175
	pesos_i(4309) := b"0000000000000000_0000000000000000_0000110111111110_0011001110100000"; -- 0.05466005951166153
	pesos_i(4310) := b"0000000000000000_0000000000000000_0011000000000001_1011111100000000"; -- 0.1875266432762146
	pesos_i(4311) := b"1111111111111111_1111111111111111_1100010101101000_1000100000000000"; -- -0.22887372970581055
	pesos_i(4312) := b"0000000000000000_0000000000000000_0000011000100111_0011100000101000"; -- 0.024035939946770668
	pesos_i(4313) := b"0000000000000000_0000000000000000_0011000111000111_1111111011000000"; -- 0.19445793330669403
	pesos_i(4314) := b"1111111111111111_1111111111111111_1100111000100101_0110110101000000"; -- -0.1947414129972458
	pesos_i(4315) := b"0000000000000000_0000000000000000_0011011110100111_1111110101000000"; -- 0.21740706264972687
	pesos_i(4316) := b"1111111111111111_1111111111111111_1100000101001100_1010010111000000"; -- -0.24492420256137848
	pesos_i(4317) := b"1111111111111111_1111111111111111_1101011001101000_1100001100000000"; -- -0.1624639630317688
	pesos_i(4318) := b"0000000000000000_0000000000000000_0000001101011111_1111100100000000"; -- 0.013183176517486572
	pesos_i(4319) := b"0000000000000000_0000000000000000_0011011011100110_1001100100000000"; -- 0.21445614099502563
	pesos_i(4320) := b"0000000000000000_0000000000000000_0100100010010011_0000110000000000"; -- 0.2834937572479248
	pesos_i(4321) := b"1111111111111111_1111111111111111_1101001010101111_1110000011000000"; -- -0.17700381577014923
	pesos_i(4322) := b"0000000000000000_0000000000000000_0011011101101110_1000100101000000"; -- 0.21653039753437042
	pesos_i(4323) := b"1111111111111111_1111111111111111_1010100100010010_1101100000000000"; -- -0.3395562171936035
	pesos_i(4324) := b"0000000000000000_0000000000000000_0000000100010110_1011011111100110"; -- 0.004252904560416937
	pesos_i(4325) := b"0000000000000000_0000000000000000_0001010111000010_1111000001100000"; -- 0.08500578254461288
	pesos_i(4326) := b"0000000000000000_0000000000000000_0000111101000011_0001001011110000"; -- 0.059617217630147934
	pesos_i(4327) := b"1111111111111111_1111111111111111_1110101001001011_1000011100000000"; -- -0.08478504419326782
	pesos_i(4328) := b"0000000000000000_0000000000000000_0001000010100111_0100001011100000"; -- 0.06505220383405685
	pesos_i(4329) := b"0000000000000000_0000000000000000_0001100011010011_0101010001000000"; -- 0.09697462618350983
	pesos_i(4330) := b"1111111111111111_1111111111111111_0111100100010111_1001111000000000"; -- -0.526983380317688
	pesos_i(4331) := b"1111111111111111_1111111111111111_1111000010111101_0010101000000000"; -- -0.059613585472106934
	pesos_i(4332) := b"0000000000000000_0000000000000000_0100111001001101_1000110100000000"; -- 0.30587083101272583
	pesos_i(4333) := b"1111111111111111_1111111111111111_1011010011110010_1010001110000000"; -- -0.2931726276874542
	pesos_i(4334) := b"0000000000000000_0000000000000000_0011101000111111_1010000101000000"; -- 0.22753341495990753
	pesos_i(4335) := b"1111111111111111_1111111111111111_0101011011011111_1010001100000000"; -- -0.6606500744819641
	pesos_i(4336) := b"0000000000000000_0000000000000000_0000010011010010_1000001011111000"; -- 0.018837152048945427
	pesos_i(4337) := b"0000000000000000_0000000000000000_0001011101100001_1110010110100000"; -- 0.09133753925561905
	pesos_i(4338) := b"0000000000000000_0000000000000000_0001000000111101_0010111000100000"; -- 0.06343353539705276
	pesos_i(4339) := b"0000000000000000_0000000000000000_0001100100001010_0110100101000000"; -- 0.09781511127948761
	pesos_i(4340) := b"1111111111111111_1111111111111111_1111011100001010_0000000110000000"; -- -0.03500357270240784
	pesos_i(4341) := b"0000000000000000_0000000000000000_0000111000010011_0111101111100000"; -- 0.05498480051755905
	pesos_i(4342) := b"0000000000000000_0000000000000000_0010010000111000_0111100100000000"; -- 0.14148670434951782
	pesos_i(4343) := b"0000000000000000_0000000000000000_0001101001111011_1001100011000000"; -- 0.10344843566417694
	pesos_i(4344) := b"1111111111111111_1111111111111111_1110101001111011_0110111000100000"; -- -0.08405410498380661
	pesos_i(4345) := b"0000000000000000_0000000000000000_0001001111011010_1100110010100000"; -- 0.07755736261606216
	pesos_i(4346) := b"1111111111111111_1111111111111111_1011111010111101_1011100010000000"; -- -0.25491759181022644
	pesos_i(4347) := b"0000000000000000_0000000000000000_0010110011100111_0000101101000000"; -- 0.17540045082569122
	pesos_i(4348) := b"1111111111111111_1111111111111111_1110101111100010_0110100111000000"; -- -0.07857646048069
	pesos_i(4349) := b"0000000000000000_0000000000000000_0000011101111110_0010001100100000"; -- 0.029268451035022736
	pesos_i(4350) := b"1111111111111111_1111111111111111_1110011000001101_0010010001100000"; -- -0.1013619676232338
	pesos_i(4351) := b"0000000000000000_0000000000000000_0001100100100011_1001000101100000"; -- 0.09819897264242172
	pesos_i(4352) := b"1111111111111111_1111111111111111_1100000001001010_1001001101000000"; -- -0.24886207282543182
	pesos_i(4353) := b"1111111111111111_1111111111111111_1101011011000001_0101010011000000"; -- -0.16111250221729279
	pesos_i(4354) := b"0000000000000000_0000000000000000_0100010111010111_1000111000000000"; -- 0.2728203535079956
	pesos_i(4355) := b"0000000000000000_0000000000000000_0010010001101000_0101110111000000"; -- 0.1422175019979477
	pesos_i(4356) := b"1111111111111111_1111111111111111_1110011100000011_0011000101100000"; -- -0.09760753065347672
	pesos_i(4357) := b"0000000000000000_0000000000000000_0011111110111011_1111010101000000"; -- 0.24896176159381866
	pesos_i(4358) := b"0000000000000000_0000000000000000_0001111100000100_0010111011100000"; -- 0.12115757912397385
	pesos_i(4359) := b"0000000000000000_0000000000000000_0011000100000110_1011011000000000"; -- 0.19150865077972412
	pesos_i(4360) := b"1111111111111111_1111111111111111_1011100011110001_0000000110000000"; -- -0.27757254242897034
	pesos_i(4361) := b"1111111111111111_1111111111111111_1100100001111110_1111100100000000"; -- -0.21681255102157593
	pesos_i(4362) := b"1111111111111111_1111111111111111_1101100000000110_0110111000000000"; -- -0.1561518907546997
	pesos_i(4363) := b"1111111111111111_1111111111111111_1110111101001101_1011111001000000"; -- -0.06521998345851898
	pesos_i(4364) := b"0000000000000000_0000000000000000_0111010111011010_1010111010000000"; -- 0.4603680670261383
	pesos_i(4365) := b"0000000000000000_0000000000000000_0111011011110011_1111111100000000"; -- 0.4646605849266052
	pesos_i(4366) := b"0000000000000000_0000000000000000_0111111110011101_0100100010000000"; -- 0.4984937012195587
	pesos_i(4367) := b"0000000000000000_0000000000000000_0011010011010001_1001000101000000"; -- 0.20632274448871613
	pesos_i(4368) := b"0000000000000000_0000000000000000_0100001100000111_0100101100000000"; -- 0.26183003187179565
	pesos_i(4369) := b"0000000000000000_0000000000000000_0000000110011000_0001101001011000"; -- 0.006227156147360802
	pesos_i(4370) := b"0000000000000000_0000000000000000_0000000100001010_1110111101111110"; -- 0.004073112737387419
	pesos_i(4371) := b"0000000000000000_0000000000000000_0000111111101110_1010011100010000"; -- 0.06223529949784279
	pesos_i(4372) := b"0000000000000000_0000000000000000_0011011111011000_0110011111000000"; -- 0.21814583241939545
	pesos_i(4373) := b"1111111111111111_1111111111111111_1110011000101101_0100001000100000"; -- -0.10087191313505173
	pesos_i(4374) := b"0000000000000000_0000000000000000_0110110010101100_0110101110000000"; -- 0.42450591921806335
	pesos_i(4375) := b"0000000000000000_0000000000000000_0001110010011111_1001100011000000"; -- 0.11181025207042694
	pesos_i(4376) := b"0000000000000000_0000000000000000_0100011101101000_1010101000000000"; -- 0.2789407968521118
	pesos_i(4377) := b"0000000000000000_0000000000000000_0111010001010010_0000011100000000"; -- 0.4543766379356384
	pesos_i(4378) := b"1111111111111111_1111111111111111_1000110011100000_0100111110000000"; -- -0.44970229268074036
	pesos_i(4379) := b"0000000000000000_0000000000000000_0001001010010001_1110110110000000"; -- 0.07253918051719666
	pesos_i(4380) := b"0000000000000000_0000000000000000_0100000110010110_0100110100000000"; -- 0.2561996579170227
	pesos_i(4381) := b"0000000000000000_0000000000000000_0110011010001010_1001011000000000"; -- 0.4005521535873413
	pesos_i(4382) := b"1111111111111111_1111111111111111_1010001101001111_0101110100000000"; -- -0.3620702624320984
	pesos_i(4383) := b"0000000000000000_0000000000000000_0001100100010001_0001101011100000"; -- 0.09791725128889084
	pesos_i(4384) := b"0000000000000000_0000000000000000_0100111101000000_1010010100000000"; -- 0.30958014726638794
	pesos_i(4385) := b"0000000000000000_0000000000000000_0011010001011100_1110110011000000"; -- 0.20454291999340057
	pesos_i(4386) := b"0000000000000000_0000000000000000_0011010100101010_1100011101000000"; -- 0.2076839953660965
	pesos_i(4387) := b"0000000000000000_0000000000000000_0101001111110100_1101100110000000"; -- 0.32795485854148865
	pesos_i(4388) := b"1111111111111111_1111111111111111_1010110010001100_1100011110000000"; -- -0.3259768784046173
	pesos_i(4389) := b"1111111111111111_1111111111111111_1011110001100011_0111011100000000"; -- -0.26410728693008423
	pesos_i(4390) := b"1111111111111111_1111111111111111_1010100111110111_0100010110000000"; -- -0.3360706865787506
	pesos_i(4391) := b"0000000000000000_0000000000000000_0110010110011110_1011010000000000"; -- 0.39695286750793457
	pesos_i(4392) := b"1111111111111111_1111111111111111_1111111010111001_1001011101110010"; -- -0.0049805971793830395
	pesos_i(4393) := b"1111111111111111_1111111111111111_1111010011100111_0010111100000000"; -- -0.04334741830825806
	pesos_i(4394) := b"0000000000000000_0000000000000000_0001110001111110_1111011111100000"; -- 0.1113123819231987
	pesos_i(4395) := b"1111111111111111_1111111111111111_1111100100000010_1110101101011000"; -- -0.02729920484125614
	pesos_i(4396) := b"1111111111111111_1111111111111111_1110010011110000_0110101110100000"; -- -0.10570647567510605
	pesos_i(4397) := b"1111111111111111_1111111111111111_1111001011000000_1111010001100000"; -- -0.051743246614933014
	pesos_i(4398) := b"0000000000000000_0000000000000000_0010101010011010_0111111110000000"; -- 0.16641995310783386
	pesos_i(4399) := b"1111111111111111_1111111111111111_1101000001111100_0000001000000000"; -- -0.18560779094696045
	pesos_i(4400) := b"1111111111111111_1111111111111111_1100000110011101_0101101110000000"; -- -0.24369266629219055
	pesos_i(4401) := b"1111111111111111_1111111111111111_1101000000000111_1000010011000000"; -- -0.18738527595996857
	pesos_i(4402) := b"0000000000000000_0000000000000000_0000101101000000_1010111110110000"; -- 0.043955784291028976
	pesos_i(4403) := b"1111111111111111_1111111111111111_1101100110010110_1001001101000000"; -- -0.15004615485668182
	pesos_i(4404) := b"0000000000000000_0000000000000000_0011110100100100_0011100000000000"; -- 0.23883390426635742
	pesos_i(4405) := b"0000000000000000_0000000000000000_0000101100100110_1101001100100000"; -- 0.043561168015003204
	pesos_i(4406) := b"1111111111111111_1111111111111111_1100000000001001_0000101010000000"; -- -0.24986204504966736
	pesos_i(4407) := b"1111111111111111_1111111111111111_1110100111101101_1100111011000000"; -- -0.08621509373188019
	pesos_i(4408) := b"1111111111111111_1111111111111111_1110110101110001_1101110100000000"; -- -0.07248133420944214
	pesos_i(4409) := b"1111111111111111_1111111111111111_0110101001101000_1100111100000000"; -- -0.5843382477760315
	pesos_i(4410) := b"0000000000000000_0000000000000000_0011010110100110_1010101010000000"; -- 0.2095743715763092
	pesos_i(4411) := b"1111111111111111_1111111111111111_1100001110111110_1001101011000000"; -- -0.235372856259346
	pesos_i(4412) := b"1111111111111111_1111111111111111_1110011011111110_0111011001100000"; -- -0.09767971187829971
	pesos_i(4413) := b"0000000000000000_0000000000000000_0111100010010010_0100001000000000"; -- 0.4709817171096802
	pesos_i(4414) := b"1111111111111111_1111111111111111_1100001001010000_1000011011000000"; -- -0.24095876514911652
	pesos_i(4415) := b"0000000000000000_0000000000000000_0000110001101111_0011011110110000"; -- 0.04857204481959343
	pesos_i(4416) := b"0000000000000000_0000000000000000_0001100111011010_0011110110000000"; -- 0.10098633170127869
	pesos_i(4417) := b"1111111111111111_1111111111111111_1100111011100000_0110100001000000"; -- -0.19188831746578217
	pesos_i(4418) := b"1111111111111111_1111111111111111_1000110001110011_0100011100000000"; -- -0.45136600732803345
	pesos_i(4419) := b"1111111111111111_1111111111111111_1110111111001011_0100000111100000"; -- -0.06330478936433792
	pesos_i(4420) := b"1111111111111111_1111111111111111_1110111011010010_0101011011000000"; -- -0.06710298359394073
	pesos_i(4421) := b"1111111111111111_1111111111111111_1110010110111011_0110000101100000"; -- -0.1026095524430275
	pesos_i(4422) := b"1111111111111111_1111111111111111_1101001100011001_0111101111000000"; -- -0.17539240419864655
	pesos_i(4423) := b"1111111111111111_1111111111111111_1100110111001000_0101100010000000"; -- -0.19616171717643738
	pesos_i(4424) := b"0000000000000000_0000000000000000_0101010010001100_1000010100000000"; -- 0.3302691578865051
	pesos_i(4425) := b"0000000000000000_0000000000000000_0000111011101011_0111101000110000"; -- 0.05828059837222099
	pesos_i(4426) := b"0000000000000000_0000000000000000_0010110111000101_0011010010000000"; -- 0.1787903606891632
	pesos_i(4427) := b"0000000000000000_0000000000000000_0010010000100010_1000001111000000"; -- 0.14115165174007416
	pesos_i(4428) := b"1111111111111111_1111111111111111_1011001100110011_1011100000000000"; -- -0.29999208450317383
	pesos_i(4429) := b"0000000000000000_0000000000000000_0101010001111000_0011011010000000"; -- 0.32995930314064026
	pesos_i(4430) := b"1111111111111111_1111111111111111_1000111011111001_1100111110000000"; -- -0.4415006935596466
	pesos_i(4431) := b"1111111111111111_1111111111111111_0111011110110001_0010011100000000"; -- -0.5324531197547913
	pesos_i(4432) := b"0000000000000000_0000000000000000_0100000111111111_1001001000000000"; -- 0.2578059434890747
	pesos_i(4433) := b"1111111111111111_1111111111111111_1001000100001100_0101101000000000"; -- -0.4334052801132202
	pesos_i(4434) := b"1111111111111111_1111111111111111_1110101011001110_0100110110100000"; -- -0.08278956264257431
	pesos_i(4435) := b"0000000000000000_0000000000000000_0110100011101011_0001010110000000"; -- 0.40983709692955017
	pesos_i(4436) := b"1111111111111111_1111111111111111_1000111110000000_0110001100000000"; -- -0.43944722414016724
	pesos_i(4437) := b"0000000000000000_0000000000000000_0000101000010101_0011011010010000"; -- 0.03938618674874306
	pesos_i(4438) := b"0000000000000000_0000000000000000_0101111011110110_1010101000000000"; -- 0.3709512948989868
	pesos_i(4439) := b"1111111111111111_1111111111111111_1001101010000100_1000101000000000"; -- -0.396415114402771
	pesos_i(4440) := b"0000000000000000_0000000000000000_0011001111100001_0010100110000000"; -- 0.20265445113182068
	pesos_i(4441) := b"0000000000000000_0000000000000000_0100010011010111_0001100110000000"; -- 0.2689071595668793
	pesos_i(4442) := b"0000000000000000_0000000000000000_0011100111100010_0010101010000000"; -- 0.22610726952552795
	pesos_i(4443) := b"0000000000000000_0000000000000000_0010110011001111_0001100110000000"; -- 0.17503508925437927
	pesos_i(4444) := b"1111111111111111_1111111111111111_1110101011100111_1101010110100000"; -- -0.08239998668432236
	pesos_i(4445) := b"1111111111111111_1111111111111111_1111001000100111_1011100101110000"; -- -0.054081354290246964
	pesos_i(4446) := b"0000000000000000_0000000000000000_0011110101000011_1001110001000000"; -- 0.23931290209293365
	pesos_i(4447) := b"0000000000000000_0000000000000000_0011101111111100_1000100111000000"; -- 0.2343221753835678
	pesos_i(4448) := b"1111111111111111_1111111111111111_1111011100101001_0100111010000000"; -- -0.03452596068382263
	pesos_i(4449) := b"1111111111111111_1111111111111111_1101101000110010_0101111000000000"; -- -0.1476689577102661
	pesos_i(4450) := b"0000000000000000_0000000000000000_0011001000111010_0010100001000000"; -- 0.1961999088525772
	pesos_i(4451) := b"1111111111111111_1111111111111111_1000110100001000_1111010110000000"; -- -0.44908204674720764
	pesos_i(4452) := b"1111111111111111_1111111111111111_1110100100010000_1010101001000000"; -- -0.08958946168422699
	pesos_i(4453) := b"1111111111111111_1111111111111111_1111001101001111_0101110110110000"; -- -0.049570221453905106
	pesos_i(4454) := b"1111111111111111_1111111111111111_1101110011100001_0110000000000000"; -- -0.13718605041503906
	pesos_i(4455) := b"1111111111111111_1111111111111111_1110000110000001_0010110001100000"; -- -0.11912272125482559
	pesos_i(4456) := b"0000000000000000_0000000000000000_0011010000000100_1000111111000000"; -- 0.20319460332393646
	pesos_i(4457) := b"0000000000000000_0000000000000000_0000101010011110_1000001011110000"; -- 0.04148119315505028
	pesos_i(4458) := b"0000000000000000_0000000000000000_0100001100010010_1100001110000000"; -- 0.2620050609111786
	pesos_i(4459) := b"0000000000000000_0000000000000000_0011100011110000_1001110001000000"; -- 0.22242142260074615
	pesos_i(4460) := b"0000000000000000_0000000000000000_0101110110000110_1101111100000000"; -- 0.3653392195701599
	pesos_i(4461) := b"1111111111111111_1111111111111111_1110001101000011_0010001000000000"; -- -0.11225688457489014
	pesos_i(4462) := b"0000000000000000_0000000000000000_0100101111100011_0110001100000000"; -- 0.29643839597702026
	pesos_i(4463) := b"1111111111111111_1111111111111111_1010001111011010_1100000010000000"; -- -0.35994336009025574
	pesos_i(4464) := b"1111111111111111_1111111111111111_1100101111000111_0011111110000000"; -- -0.20399096608161926
	pesos_i(4465) := b"0000000000000000_0000000000000000_0011000001100100_1010110001000000"; -- 0.18903614580631256
	pesos_i(4466) := b"0000000000000000_0000000000000000_0100010111101110_1100100010000000"; -- 0.27317479252815247
	pesos_i(4467) := b"0000000000000000_0000000000000000_0101111100111001_1000110010000000"; -- 0.37197187542915344
	pesos_i(4468) := b"1111111111111111_1111111111111111_1110101000001111_0001011011100000"; -- -0.08570725470781326
	pesos_i(4469) := b"0000000000000000_0000000000000000_0100111000101100_0011001000000000"; -- 0.30536186695098877
	pesos_i(4470) := b"0000000000000000_0000000000000000_0111000001101100_1101001110000000"; -- 0.43916055560112
	pesos_i(4471) := b"1111111111111111_1111111111111111_1000000001001110_0000110000000000"; -- -0.4988090991973877
	pesos_i(4472) := b"0000000000000000_0000000000000000_0100111110010101_1111111100000000"; -- 0.3108825087547302
	pesos_i(4473) := b"0000000000000000_0000000000000000_0101110100100111_1101100110000000"; -- 0.36388930678367615
	pesos_i(4474) := b"0000000000000000_0000000000000000_0001101000011110_1101100010100000"; -- 0.10203317552804947
	pesos_i(4475) := b"0000000000000000_0000000000000000_0010010100001011_0101111010000000"; -- 0.14470472931861877
	pesos_i(4476) := b"0000000000000000_0000000000000000_0101000100010010_0110000100000000"; -- 0.3166866898536682
	pesos_i(4477) := b"0000000000000000_0000000000000000_0001111110100000_1001000000100000"; -- 0.12354374676942825
	pesos_i(4478) := b"0000000000000000_0000000000000000_0010100111111101_1011111100000000"; -- 0.1640281081199646
	pesos_i(4479) := b"0000000000000000_0000000000000000_0010100101101011_0000000110000000"; -- 0.16178902983665466
	pesos_i(4480) := b"0000000000000000_0000000000000000_1101000001010101_1101100100000000"; -- 0.8138099312782288
	pesos_i(4481) := b"0000000000000000_0000000000000000_0001101111010101_0010011010100000"; -- 0.10872117429971695
	pesos_i(4482) := b"1111111111111111_1111111111111111_1100000101101110_1111100000000000"; -- -0.2444005012512207
	pesos_i(4483) := b"1111111111111111_1111111111111111_1111110001011111_0110111101100000"; -- -0.014168776571750641
	pesos_i(4484) := b"0000000000000000_0000000000000000_0111011010110011_0001001000000000"; -- 0.46366989612579346
	pesos_i(4485) := b"0000000000000000_0000000000000000_0111001100111110_1110111010000000"; -- 0.45017901062965393
	pesos_i(4486) := b"0000000000000000_0000000000000000_0100100011011000_0100000110000000"; -- 0.2845498025417328
	pesos_i(4487) := b"1111111111111111_1111111111111111_0110001000010110_1100001000000000"; -- -0.6168402433395386
	pesos_i(4488) := b"0000000000000000_0000000000000000_0000010000011000_0011011111000000"; -- 0.015994533896446228
	pesos_i(4489) := b"0000000000000000_0000000000000000_0110101011000010_0000010110000000"; -- 0.41702303290367126
	pesos_i(4490) := b"1111111111111111_1111111111111111_1101110000011101_0001101110000000"; -- -0.14018085598945618
	pesos_i(4491) := b"1111111111111111_1111111111111111_1011100001110010_1011010110000000"; -- -0.27949967980384827
	pesos_i(4492) := b"1111111111111111_1111111111111111_1100011101010001_1010110101000000"; -- -0.22140996158123016
	pesos_i(4493) := b"0000000000000000_0000000000000000_0010010011110100_1000001001000000"; -- 0.144355908036232
	pesos_i(4494) := b"0000000000000000_0000000000000000_0000001100010001_0010110001110000"; -- 0.011980798095464706
	pesos_i(4495) := b"1111111111111111_1111111111111111_1001101001100011_1111101110000000"; -- -0.3969118893146515
	pesos_i(4496) := b"0000000000000000_0000000000000000_0010111000110101_1011100100000000"; -- 0.18050724267959595
	pesos_i(4497) := b"0000000000000000_0000000000000000_1000110001100110_0111000000000000"; -- 0.5484380722045898
	pesos_i(4498) := b"0000000000000000_0000000000000000_0111000100111101_1011011110000000"; -- 0.4423479735851288
	pesos_i(4499) := b"0000000000000000_0000000000000000_0100100110100111_0011011110000000"; -- 0.28770777583122253
	pesos_i(4500) := b"0000000000000000_0000000000000000_0110010101110010_0110101100000000"; -- 0.39627712965011597
	pesos_i(4501) := b"0000000000000000_0000000000000000_0011011110110001_0101111011000000"; -- 0.21755020320415497
	pesos_i(4502) := b"1111111111111111_1111111111111111_1010110001100111_1111010010000000"; -- -0.3265387713909149
	pesos_i(4503) := b"0000000000000000_0000000000000000_0101010101001100_0011011000000000"; -- 0.33319413661956787
	pesos_i(4504) := b"0000000000000000_0000000000000000_0101010101101101_1011000010000000"; -- 0.33370497822761536
	pesos_i(4505) := b"1111111111111111_1111111111111111_1111000101110001_1110010110110000"; -- -0.05685581639409065
	pesos_i(4506) := b"0000000000000000_0000000000000000_0001100110000110_0111100001000000"; -- 0.09970809519290924
	pesos_i(4507) := b"0000000000000000_0000000000000000_0011000000110001_0100100111000000"; -- 0.18825207650661469
	pesos_i(4508) := b"1111111111111111_1111111111111111_1001011010000001_0111110010000000"; -- -0.41208669543266296
	pesos_i(4509) := b"0000000000000000_0000000000000000_0010111110100001_1000010011000000"; -- 0.18605832755565643
	pesos_i(4510) := b"1111111111111111_1111111111111111_1011100000111000_1111001000000000"; -- -0.28038108348846436
	pesos_i(4511) := b"1111111111111111_1111111111111111_1101111010001111_0011110000000000"; -- -0.13062691688537598
	pesos_i(4512) := b"1111111111111111_1111111111111111_1111000010011001_0001010101110000"; -- -0.06016412749886513
	pesos_i(4513) := b"1111111111111111_1111111111111111_1110011011110100_1001100010000000"; -- -0.09783026576042175
	pesos_i(4514) := b"0000000000000000_0000000000000000_0010100100011100_0010111111000000"; -- 0.16058634221553802
	pesos_i(4515) := b"1111111111111111_1111111111111111_1001111100001010_1101000110000000"; -- -0.37874117493629456
	pesos_i(4516) := b"1111111111111111_1111111111111111_1110101000100100_0000100001100000"; -- -0.08538768440485
	pesos_i(4517) := b"0000000000000000_0000000000000000_1010010010111111_1011111100000000"; -- 0.6435508131980896
	pesos_i(4518) := b"0000000000000000_0000000000000000_0000111100010100_1101001011010000"; -- 0.05891149118542671
	pesos_i(4519) := b"1111111111111111_1111111111111111_1001000001010101_0100110100000000"; -- -0.4361984133720398
	pesos_i(4520) := b"0000000000000000_0000000000000000_0001011101010001_1001011111100000"; -- 0.09108876436948776
	pesos_i(4521) := b"0000000000000000_0000000000000000_0010110001010110_1100110110000000"; -- 0.17319950461387634
	pesos_i(4522) := b"1111111111111111_1111111111111111_1111101011100010_1101011000011000"; -- -0.01997625268995762
	pesos_i(4523) := b"1111111111111111_1111111111111111_1101111101101101_1010111011000000"; -- -0.127232626080513
	pesos_i(4524) := b"1111111111111111_1111111111111111_1101000100101011_0100101000000000"; -- -0.18293321132659912
	pesos_i(4525) := b"0000000000000000_0000000000000000_0011111010000000_1010011010000000"; -- 0.2441505491733551
	pesos_i(4526) := b"1111111111111111_1111111111111111_1110110100111100_0111000110000000"; -- -0.073296457529068
	pesos_i(4527) := b"1111111111111111_1111111111111111_1111111111011001_1001001110100001"; -- -0.0005862934631295502
	pesos_i(4528) := b"0000000000000000_0000000000000000_0101101010000010_0100001000000000"; -- 0.3535500764846802
	pesos_i(4529) := b"0000000000000000_0000000000000000_0110110111110001_0001111100000000"; -- 0.42946046590805054
	pesos_i(4530) := b"0000000000000000_0000000000000000_1000001000110010_0010001000000000"; -- 0.5085774660110474
	pesos_i(4531) := b"1111111111111111_1111111111111111_1110101100101011_1010000101100000"; -- -0.08136550337076187
	pesos_i(4532) := b"1111111111111111_1111111111111111_1111011001101101_0101010011100000"; -- -0.03739423304796219
	pesos_i(4533) := b"0000000000000000_0000000000000000_0100010010001010_0000111110000000"; -- 0.267731636762619
	pesos_i(4534) := b"0000000000000000_0000000000000000_1000110100011100_1010011100000000"; -- 0.5512184500694275
	pesos_i(4535) := b"1111111111111111_1111111111111111_1111110001010010_0011010000111100"; -- -0.01437066588550806
	pesos_i(4536) := b"0000000000000000_0000000000000000_0010001111111111_1011000011000000"; -- 0.14062027633190155
	pesos_i(4537) := b"1111111111111111_1111111111111111_1010000111010011_0100011000000000"; -- -0.3678699731826782
	pesos_i(4538) := b"1111111111111111_1111111111111111_1110110000010011_0110101111100000"; -- -0.07782865315675735
	pesos_i(4539) := b"1111111111111111_1111111111111111_1111100110100000_1001011010100000"; -- -0.024893365800380707
	pesos_i(4540) := b"0000000000000000_0000000000000000_0011100011011000_1100100010000000"; -- 0.22205784916877747
	pesos_i(4541) := b"0000000000000000_0000000000000000_0111100001010101_0101010000000000"; -- 0.47005200386047363
	pesos_i(4542) := b"1111111111111111_1111111111111111_1011111110110011_0110100010000000"; -- -0.25116869807243347
	pesos_i(4543) := b"0000000000000000_0000000000000000_0011101000001011_1111100001000000"; -- 0.226745143532753
	pesos_i(4544) := b"0000000000000000_0000000000000000_0100101010101011_1001100100000000"; -- 0.29168087244033813
	pesos_i(4545) := b"1111111111111111_1111111111111111_1100111111001111_0001001010000000"; -- -0.18824657797813416
	pesos_i(4546) := b"0000000000000000_0000000000000000_0111010100011010_0001011110000000"; -- 0.4574293792247772
	pesos_i(4547) := b"0000000000000000_0000000000000000_0010100101001101_0011101001000000"; -- 0.16133464872837067
	pesos_i(4548) := b"1111111111111111_1111111111111111_1101100100110111_1111111011000000"; -- -0.15148933231830597
	pesos_i(4549) := b"0000000000000000_0000000000000000_1000010011101000_0010110000000000"; -- 0.5191676616668701
	pesos_i(4550) := b"0000000000000000_0000000000000000_0011100111011011_0000011100000000"; -- 0.22599834203720093
	pesos_i(4551) := b"0000000000000000_0000000000000000_0010010010110100_1001101110000000"; -- 0.14338085055351257
	pesos_i(4552) := b"1111111111111111_1111111111111111_1010100000110011_0001000000000000"; -- -0.3429708480834961
	pesos_i(4553) := b"1111111111111111_1111111111111111_0110010000100000_1101111100000000"; -- -0.6088734269142151
	pesos_i(4554) := b"0000000000000000_0000000000000000_0011011011101101_0110001011000000"; -- 0.21455971896648407
	pesos_i(4555) := b"0000000000000000_0000000000000000_0100101000100010_0001100100000000"; -- 0.2895827889442444
	pesos_i(4556) := b"0000000000000000_0000000000000000_0100100111111010_0011011000000000"; -- 0.28897416591644287
	pesos_i(4557) := b"0000000000000000_0000000000000000_0010000000000010_0101011000000000"; -- 0.12503564357757568
	pesos_i(4558) := b"1111111111111111_1111111111111111_1100110001101010_1011001000000000"; -- -0.20149695873260498
	pesos_i(4559) := b"0000000000000000_0000000000000000_0100100010001100_0000010110000000"; -- 0.28338655829429626
	pesos_i(4560) := b"1111111111111111_1111111111111111_1111000001111101_0100010110010000"; -- -0.06058850511908531
	pesos_i(4561) := b"1111111111111111_1111111111111111_1001101000010110_0110010100000000"; -- -0.3980957865715027
	pesos_i(4562) := b"0000000000000000_0000000000000000_0101101111111100_0101011000000000"; -- 0.3593190908432007
	pesos_i(4563) := b"0000000000000000_0000000000000000_0101100010000100_0101001110000000"; -- 0.34576913714408875
	pesos_i(4564) := b"0000000000000000_0000000000000000_0001011110101111_0100001100100000"; -- 0.09251803904771805
	pesos_i(4565) := b"1111111111111111_1111111111111111_1110101010011100_0011000110000000"; -- -0.08355417847633362
	pesos_i(4566) := b"1111111111111111_1111111111111111_1010101101110010_1000101100000000"; -- -0.3302834630012512
	pesos_i(4567) := b"1111111111111111_1111111111111110_1100111101100110_1101010000000000"; -- -1.1898372173309326
	pesos_i(4568) := b"1111111111111111_1111111111111111_1011111011110101_1101001100000000"; -- -0.2540615200996399
	pesos_i(4569) := b"0000000000000000_0000000000000000_0000110001100101_1000110000000000"; -- 0.048424482345581055
	pesos_i(4570) := b"0000000000000000_0000000000000000_1000001011010101_1111100100000000"; -- 0.5110774636268616
	pesos_i(4571) := b"1111111111111111_1111111111111111_1111010001001100_0001100000110000"; -- -0.045713890343904495
	pesos_i(4572) := b"1111111111111111_1111111111111111_1110001011101011_1010010011100000"; -- -0.11359185725450516
	pesos_i(4573) := b"0000000000000000_0000000000000000_0011011011111100_0101110111000000"; -- 0.2147883027791977
	pesos_i(4574) := b"0000000000000000_0000000000000000_0101100100011011_1011000000000000"; -- 0.34807872772216797
	pesos_i(4575) := b"0000000000000000_0000000000000000_0011111101011110_1101110100000000"; -- 0.24754124879837036
	pesos_i(4576) := b"0000000000000000_0000000000000000_0010011100010110_1110000000000000"; -- 0.1526927947998047
	pesos_i(4577) := b"1111111111111111_1111111111111111_1100011111010010_0010100000000000"; -- -0.21944952011108398
	pesos_i(4578) := b"1111111111111111_1111111111111111_1000010010110001_0011110100000000"; -- -0.4816705584526062
	pesos_i(4579) := b"0000000000000000_0000000000000000_0001011111011011_0001111001000000"; -- 0.09318722784519196
	pesos_i(4580) := b"1111111111111111_1111111111111111_1110100010000010_1001111000000000"; -- -0.09175693988800049
	pesos_i(4581) := b"1111111111111111_1111111111111111_1101100111001100_0000101000000000"; -- -0.14923036098480225
	pesos_i(4582) := b"1111111111111111_1111111111111111_1111000000110011_1100010110000000"; -- -0.06171002984046936
	pesos_i(4583) := b"0000000000000000_0000000000000000_0010010010000001_1110000011000000"; -- 0.14260677993297577
	pesos_i(4584) := b"0000000000000000_0000000000000000_1000101100110011_1111100100000000"; -- 0.5437617897987366
	pesos_i(4585) := b"0000000000000000_0000000000000000_0001100010110001_0001000101000000"; -- 0.09645183384418488
	pesos_i(4586) := b"0000000000000000_0000000000000000_0001010000101001_0011011011100000"; -- 0.07875388115644455
	pesos_i(4587) := b"1111111111111111_1111111111111111_1110110000011000_0110010111100000"; -- -0.07775271683931351
	pesos_i(4588) := b"0000000000000000_0000000000000000_1000100111010100_1011111100000000"; -- 0.5384024977684021
	pesos_i(4589) := b"0000000000000000_0000000000000000_0000000011111110_1100110000001010"; -- 0.0038878940977156162
	pesos_i(4590) := b"1111111111111111_1111111111111111_1100000010000010_0111001000000000"; -- -0.2480095624923706
	pesos_i(4591) := b"1111111111111111_1111111111111111_1100011101010000_0000100010000000"; -- -0.2214350402355194
	pesos_i(4592) := b"0000000000000000_0000000000000000_0110100011101100_1111001110000000"; -- 0.4098655879497528
	pesos_i(4593) := b"0000000000000000_0000000000000000_1001110111001001_1101101000000000"; -- 0.6163612604141235
	pesos_i(4594) := b"0000000000000000_0000000000000000_0111100001101001_0000100100000000"; -- 0.4703527092933655
	pesos_i(4595) := b"1111111111111111_1111111111111111_1101011010100011_1011100010000000"; -- -0.16156432032585144
	pesos_i(4596) := b"0000000000000000_0000000000000000_0010001001100001_1001010110000000"; -- 0.13430151343345642
	pesos_i(4597) := b"0000000000000000_0000000000000000_0100101101111100_0100100010000000"; -- 0.2948651611804962
	pesos_i(4598) := b"1111111111111111_1111111111111111_1100101101001010_0111001011000000"; -- -0.20589525997638702
	pesos_i(4599) := b"1111111111111111_1111111111111111_1011000111010000_1101110110000000"; -- -0.30540671944618225
	pesos_i(4600) := b"0000000000000000_0000000000000000_0100000100110001_0100001000000000"; -- 0.2546578645706177
	pesos_i(4601) := b"1111111111111111_1111111111111111_1010110111101110_0010101110000000"; -- -0.32058456540107727
	pesos_i(4602) := b"0000000000000000_0000000000000000_0110111101100101_1100111000000000"; -- 0.43514716625213623
	pesos_i(4603) := b"0000000000000000_0000000000000000_0000011011111000_1110001110100000"; -- 0.027235247194767
	pesos_i(4604) := b"1111111111111111_1111111111111111_1001010010000100_1001000110000000"; -- -0.4198521673679352
	pesos_i(4605) := b"0000000000000000_0000000000000000_0011000101110001_0011111101000000"; -- 0.19313426315784454
	pesos_i(4606) := b"0000000000000000_0000000000000001_0000011111010111_0010000000000000"; -- 1.0306262969970703
	pesos_i(4607) := b"1111111111111111_1111111111111111_1110010000100111_1111001111100000"; -- -0.1087653711438179
	pesos_i(4608) := b"0000000000000000_0000000000000000_1000011001110001_0010111100000000"; -- 0.5251645445823669
	pesos_i(4609) := b"0000000000000000_0000000000000000_0000100110001100_0010010011000000"; -- 0.037294670939445496
	pesos_i(4610) := b"1111111111111111_1111111111111111_1010000111000010_1011111110000000"; -- -0.3681221306324005
	pesos_i(4611) := b"0000000000000000_0000000000000000_0100000010110011_0011000100000000"; -- 0.2527342438697815
	pesos_i(4612) := b"0000000000000000_0000000000000000_1000011101101110_1001100100000000"; -- 0.5290313363075256
	pesos_i(4613) := b"1111111111111111_1111111111111111_1111010111111001_0011011110000000"; -- -0.039166003465652466
	pesos_i(4614) := b"1111111111111111_1111111111111111_1110110110111111_0111001111000000"; -- -0.07129742205142975
	pesos_i(4615) := b"1111111111111111_1111111111111111_1010001110011100_1011100010000000"; -- -0.36088988184928894
	pesos_i(4616) := b"0000000000000000_0000000000000000_1000001110101010_1101000000000000"; -- 0.5143251419067383
	pesos_i(4617) := b"1111111111111111_1111111111111111_1110110110000011_1101010011100000"; -- -0.07220716029405594
	pesos_i(4618) := b"0000000000000000_0000000000000000_0010011010101101_0100011011000000"; -- 0.15108148753643036
	pesos_i(4619) := b"0000000000000000_0000000000000000_0100000000100100_0101101110000000"; -- 0.25055477023124695
	pesos_i(4620) := b"1111111111111111_1111111111111111_1101101111001000_1010110110000000"; -- -0.14146915078163147
	pesos_i(4621) := b"1111111111111111_1111111111111111_1111110001110110_0100011010111100"; -- -0.013820246793329716
	pesos_i(4622) := b"1111111111111111_1111111111111111_1010000011111100_0001111110000000"; -- -0.3711529076099396
	pesos_i(4623) := b"1111111111111111_1111111111111111_1011010101001101_1100010010000000"; -- -0.29178211092948914
	pesos_i(4624) := b"0000000000000000_0000000000000000_0111000101000011_0010000100000000"; -- 0.4424305558204651
	pesos_i(4625) := b"0000000000000000_0000000000000000_0010101010001001_1101101110000000"; -- 0.1661660373210907
	pesos_i(4626) := b"1111111111111111_1111111111111111_1110010111101010_1000110111100000"; -- -0.10188973695039749
	pesos_i(4627) := b"0000000000000000_0000000000000000_0000010000110111_1101001011000000"; -- 0.016476795077323914
	pesos_i(4628) := b"0000000000000000_0000000000000000_0001111001010100_1000000000000000"; -- 0.11847686767578125
	pesos_i(4629) := b"0000000000000000_0000000000000000_1000101011111111_1010100100000000"; -- 0.5429635643959045
	pesos_i(4630) := b"1111111111111111_1111111111111111_0111011101011010_1001011100000000"; -- -0.5337739586830139
	pesos_i(4631) := b"0000000000000000_0000000000000000_0110010100011001_1101110010000000"; -- 0.3949258625507355
	pesos_i(4632) := b"0000000000000000_0000000000000000_0111001111110010_1110100110000000"; -- 0.45292529463768005
	pesos_i(4633) := b"0000000000000000_0000000000000000_0010101100110100_0011001101000000"; -- 0.16876526176929474
	pesos_i(4634) := b"0000000000000000_0000000000000000_0000001111101110_1000111001100000"; -- 0.015358828008174896
	pesos_i(4635) := b"0000000000000000_0000000000000000_0110000111011010_0001101100000000"; -- 0.38223427534103394
	pesos_i(4636) := b"1111111111111111_1111111111111111_1110010101100111_1010111111000000"; -- -0.10388661921024323
	pesos_i(4637) := b"1111111111111111_1111111111111111_1011001101111110_1010001000000000"; -- -0.2988489866256714
	pesos_i(4638) := b"0000000000000000_0000000000000000_0001010011100110_1110111011000000"; -- 0.08164875209331512
	pesos_i(4639) := b"0000000000000000_0000000000000000_0000110000000110_1110010011000000"; -- 0.04698018729686737
	pesos_i(4640) := b"0000000000000000_0000000000000000_0110001101011101_0111100000000000"; -- 0.38814496994018555
	pesos_i(4641) := b"1111111111111111_1111111111111111_1100100101110100_1101000001000000"; -- -0.21306131780147552
	pesos_i(4642) := b"1111111111111111_1111111111111111_1001110010111110_1001010110000000"; -- -0.3877169191837311
	pesos_i(4643) := b"1111111111111111_1111111111111111_1101110101000010_0101001111000000"; -- -0.13570667803287506
	pesos_i(4644) := b"1111111111111111_1111111111111111_1000110100111011_1111110110000000"; -- -0.44830337166786194
	pesos_i(4645) := b"0000000000000000_0000000000000000_0011101100101001_1000000011000000"; -- 0.23110203444957733
	pesos_i(4646) := b"0000000000000000_0000000000000000_0101000010001110_1010111010000000"; -- 0.3146771490573883
	pesos_i(4647) := b"1111111111111111_1111111111111111_0101011010011110_0011001100000000"; -- -0.6616485714912415
	pesos_i(4648) := b"1111111111111111_1111111111111111_1101001100101100_0010011001000000"; -- -0.17510758340358734
	pesos_i(4649) := b"1111111111111111_1111111111111111_1111000110010100_0100001010100000"; -- -0.05633147805929184
	pesos_i(4650) := b"1111111111111111_1111111111111111_1110010011110000_0101011011100000"; -- -0.10570771247148514
	pesos_i(4651) := b"0000000000000000_0000000000000000_0001010100011110_0111100111000000"; -- 0.0824962705373764
	pesos_i(4652) := b"0000000000000000_0000000000000000_0011110110011010_0101010101000000"; -- 0.2406361848115921
	pesos_i(4653) := b"1111111111111111_1111111111111111_1010010100110101_0100000100000000"; -- -0.3546561598777771
	pesos_i(4654) := b"0000000000000000_0000000000000000_0101010100010000_1101010110000000"; -- 0.33228811621665955
	pesos_i(4655) := b"1111111111111111_1111111111111111_1010110011001101_0010111010000000"; -- -0.32499417662620544
	pesos_i(4656) := b"1111111111111111_1111111111111111_1101100111101010_0101011110000000"; -- -0.14876797795295715
	pesos_i(4657) := b"0000000000000000_0000000000000000_0101110001101101_1001110000000000"; -- 0.36104750633239746
	pesos_i(4658) := b"0000000000000000_0000000000000000_0101010001000010_1101111000000000"; -- 0.32914531230926514
	pesos_i(4659) := b"0000000000000000_0000000000000000_0010011110001011_0010111111000000"; -- 0.15446756780147552
	pesos_i(4660) := b"1111111111111111_1111111111111111_1010010011001101_0101001110000000"; -- -0.35624197125434875
	pesos_i(4661) := b"0000000000000000_0000000000000000_0101110110111101_1010101100000000"; -- 0.3661753535270691
	pesos_i(4662) := b"1111111111111111_1111111111111111_1101111100000111_1101110001000000"; -- -0.12878631055355072
	pesos_i(4663) := b"0000000000000000_0000000000000000_0011010100100001_1110010000000000"; -- 0.2075483798980713
	pesos_i(4664) := b"0000000000000000_0000000000000000_0101001001101110_1101010100000000"; -- 0.32200366258621216
	pesos_i(4665) := b"0000000000000000_0000000000000000_0011101001111101_0101110001000000"; -- 0.22847534716129303
	pesos_i(4666) := b"0000000000000000_0000000000000000_0111100010001100_1100000010000000"; -- 0.47089770436286926
	pesos_i(4667) := b"1111111111111111_1111111111111111_1101110000010100_1101001101000000"; -- -0.1403072327375412
	pesos_i(4668) := b"0000000000000000_0000000000000000_0110100111101110_1000010100000000"; -- 0.4137957692146301
	pesos_i(4669) := b"0000000000000000_0000000000000000_0001000011011001_1111001101000000"; -- 0.06582565605640411
	pesos_i(4670) := b"0000000000000000_0000000000000000_0010010000111000_0101101100000000"; -- 0.14148491621017456
	pesos_i(4671) := b"1111111111111111_1111111111111111_1111101100010001_1011100100100000"; -- -0.019260816276073456
	pesos_i(4672) := b"0000000000000000_0000000000000000_0011111010100000_1100000011000000"; -- 0.24464039504528046
	pesos_i(4673) := b"0000000000000000_0000000000000000_0011001110111010_1110100101000000"; -- 0.20207078754901886
	pesos_i(4674) := b"0000000000000000_0000000000000000_0001111100100110_0110001101100000"; -- 0.12167950719594955
	pesos_i(4675) := b"1111111111111111_1111111111111111_1011101011011110_0011010100000000"; -- -0.2700468897819519
	pesos_i(4676) := b"0000000000000000_0000000000000000_0010110000101010_0010111101000000"; -- 0.17251868546009064
	pesos_i(4677) := b"0000000000000000_0000000000000000_0011111110000101_0111010010000000"; -- 0.24813011288642883
	pesos_i(4678) := b"0000000000000000_0000000000000000_0010000011110111_1100001100000000"; -- 0.1287805438041687
	pesos_i(4679) := b"0000000000000000_0000000000000000_1000011110100111_1110110000000000"; -- 0.5299060344696045
	pesos_i(4680) := b"1111111111111111_1111111111111111_1101100110111111_1100101110000000"; -- -0.1494171917438507
	pesos_i(4681) := b"1111111111111111_1111111111111111_1010100011101101_0100010000000000"; -- -0.3401296138763428
	pesos_i(4682) := b"0000000000000000_0000000000000000_0001110001110001_1111011111000000"; -- 0.1111140102148056
	pesos_i(4683) := b"0000000000000000_0000000000000000_0110101111010101_1100011100000000"; -- 0.4212307333946228
	pesos_i(4684) := b"0000000000000000_0000000000000000_0001101111110011_1100100101100000"; -- 0.10918863862752914
	pesos_i(4685) := b"0000000000000000_0000000000000000_0000111101011100_1110111110000000"; -- 0.060011833906173706
	pesos_i(4686) := b"0000000000000000_0000000000000000_0011011010000000_1101101001000000"; -- 0.21290363371372223
	pesos_i(4687) := b"0000000000000000_0000000000000000_0100000000010111_1011010010000000"; -- 0.25036171078681946
	pesos_i(4688) := b"0000000000000000_0000000000000000_0111101101001011_1001010100000000"; -- 0.48162204027175903
	pesos_i(4689) := b"1111111111111111_1111111111111111_1110010000011001_0101110001000000"; -- -0.10898803174495697
	pesos_i(4690) := b"0000000000000000_0000000000000000_0100000010101100_0110111000000000"; -- 0.2526310682296753
	pesos_i(4691) := b"0000000000000000_0000000000000000_0000101101011000_0111011001010000"; -- 0.04431857541203499
	pesos_i(4692) := b"0000000000000000_0000000000000000_0100111110101110_0100100010000000"; -- 0.3112531006336212
	pesos_i(4693) := b"1111111111111111_1111111111111111_1111010101100101_0001111101010000"; -- -0.04142574593424797
	pesos_i(4694) := b"1111111111111111_1111111111111111_1100101110001100_0010010000000000"; -- -0.20489287376403809
	pesos_i(4695) := b"0000000000000000_0000000000000000_0011000011001001_1000010100000000"; -- 0.19057494401931763
	pesos_i(4696) := b"1111111111111111_1111111111111111_0111011100011110_1110111100000000"; -- -0.5346842408180237
	pesos_i(4697) := b"1111111111111111_1111111111111111_1100111110110011_1011011101000000"; -- -0.1886640042066574
	pesos_i(4698) := b"0000000000000000_0000000000000000_1000101000101001_0110101000000000"; -- 0.5396944284439087
	pesos_i(4699) := b"0000000000000000_0000000000000000_0001110000110001_0000101000100000"; -- 0.11012328416109085
	pesos_i(4700) := b"0000000000000000_0000000000000000_1001101010000000_1011011100000000"; -- 0.6035265326499939
	pesos_i(4701) := b"0000000000000000_0000000000000000_0100011110100001_0111011100000000"; -- 0.27980750799179077
	pesos_i(4702) := b"0000000000000000_0000000000000000_0101001100001101_1011011010000000"; -- 0.324427992105484
	pesos_i(4703) := b"1111111111111111_1111111111111111_1111000010011000_0001111101000000"; -- -0.06017880141735077
	pesos_i(4704) := b"0000000000000000_0000000000000000_0011010011110000_1010111111000000"; -- 0.20679758489131927
	pesos_i(4705) := b"1111111111111111_1111111111111111_1100110001001010_0110011100000000"; -- -0.20198971033096313
	pesos_i(4706) := b"0000000000000000_0000000000000000_0000010010010000_1001000101100000"; -- 0.017830930650234222
	pesos_i(4707) := b"0000000000000000_0000000000000000_0001010011101110_0011110001100000"; -- 0.08176019042730331
	pesos_i(4708) := b"1111111111111111_1111111111111111_1010011011011011_0111010010000000"; -- -0.34821388125419617
	pesos_i(4709) := b"1111111111111111_1111111111111111_0100100011110110_0011011100000000"; -- -0.7149930596351624
	pesos_i(4710) := b"1111111111111111_1111111111111111_1100111001001100_1011000110000000"; -- -0.19414225220680237
	pesos_i(4711) := b"0000000000000000_0000000000000000_0001010100001000_1011010111100000"; -- 0.08216416090726852
	pesos_i(4712) := b"0000000000000000_0000000000000000_0001110000111011_0010101010100000"; -- 0.11027780920267105
	pesos_i(4713) := b"0000000000000000_0000000000000000_0100111011101010_1100010000000000"; -- 0.308269739151001
	pesos_i(4714) := b"1111111111111111_1111111111111111_1110011110110000_0101001010100000"; -- -0.09496577829122543
	pesos_i(4715) := b"1111111111111111_1111111111111111_1011111001100100_0011101100000000"; -- -0.25628310441970825
	pesos_i(4716) := b"0000000000000000_0000000000000000_0010011110100011_0111011100000000"; -- 0.15483802556991577
	pesos_i(4717) := b"0000000000000000_0000000000000000_0001100001001010_1111011110000000"; -- 0.09489390254020691
	pesos_i(4718) := b"1111111111111111_1111111111111111_1111010011101000_0001101111000000"; -- -0.04333330690860748
	pesos_i(4719) := b"1111111111111111_1111111111111111_1111010010100000_1111101011000000"; -- -0.04441864788532257
	pesos_i(4720) := b"0000000000000000_0000000000000000_0101010110101000_1010011110000000"; -- 0.3346047103404999
	pesos_i(4721) := b"0000000000000000_0000000000000000_0101000100110000_0111001000000000"; -- 0.3171454668045044
	pesos_i(4722) := b"0000000000000000_0000000000000000_0101111100001111_1100010000000000"; -- 0.3713343143463135
	pesos_i(4723) := b"0000000000000000_0000000000000000_1000001011010101_0110111000000000"; -- 0.5110691785812378
	pesos_i(4724) := b"0000000000000000_0000000000000000_0100110010111111_1010110100000000"; -- 0.29979974031448364
	pesos_i(4725) := b"0000000000000000_0000000000000000_0010100101110000_1010111100000000"; -- 0.1618756651878357
	pesos_i(4726) := b"0000000000000000_0000000000000000_0010101001010111_0010011011000000"; -- 0.16539232432842255
	pesos_i(4727) := b"0000000000000000_0000000000000000_0100011001111100_1001011110000000"; -- 0.27533861994743347
	pesos_i(4728) := b"0000000000000000_0000000000000000_0100100000111110_1000001100000000"; -- 0.2822038531303406
	pesos_i(4729) := b"1111111111111111_1111111111111111_1100001011010000_1111000011000000"; -- -0.23899932205677032
	pesos_i(4730) := b"0000000000000000_0000000000000000_0011111100000010_1100101100000000"; -- 0.2461363673210144
	pesos_i(4731) := b"0000000000000000_0000000000000000_0100111000100011_1111110010000000"; -- 0.3052366077899933
	pesos_i(4732) := b"1111111111111111_1111111111111111_1010010011011001_1001101000000000"; -- -0.3560546636581421
	pesos_i(4733) := b"0000000000000000_0000000000000000_0011100010011100_0110011011000000"; -- 0.22113649547100067
	pesos_i(4734) := b"0000000000000000_0000000000000000_0011100101100101_1001010110000000"; -- 0.22420629858970642
	pesos_i(4735) := b"1111111111111111_1111111111111111_1101110000011111_0001010100000000"; -- -0.14015072584152222
	pesos_i(4736) := b"0000000000000000_0000000000000000_0000011000100011_0011111001111000"; -- 0.023975281044840813
	pesos_i(4737) := b"0000000000000000_0000000000000000_0100011110001111_1010100010000000"; -- 0.27953580021858215
	pesos_i(4738) := b"1111111111111111_1111111111111111_1101000010101011_1110100000000000"; -- -0.1848769187927246
	pesos_i(4739) := b"0000000000000000_0000000000000000_0100001100011111_1001100100000000"; -- 0.26220089197158813
	pesos_i(4740) := b"1111111111111111_1111111111111111_1110001100011111_0001011101100000"; -- -0.11280683428049088
	pesos_i(4741) := b"1111111111111111_1111111111111111_0111010011110111_1000000000000000"; -- -0.5430984497070312
	pesos_i(4742) := b"0000000000000000_0000000000000000_0001101000100011_1010010101000000"; -- 0.10210640728473663
	pesos_i(4743) := b"0000000000000000_0000000000000000_0001010101010000_0001101000000000"; -- 0.08325350284576416
	pesos_i(4744) := b"0000000000000000_0000000000000000_0000110001011101_1101110101100000"; -- 0.04830726236104965
	pesos_i(4745) := b"1111111111111111_1111111111111111_1101010110000001_1100101001000000"; -- -0.16598831117153168
	pesos_i(4746) := b"0000000000000000_0000000000000000_0101011001010101_0111101100000000"; -- 0.3372418284416199
	pesos_i(4747) := b"0000000000000000_0000000000000000_0000100111001111_1011000011010000"; -- 0.03832535818219185
	pesos_i(4748) := b"0000000000000000_0000000000000000_0010100001110010_1101001000000000"; -- 0.15800201892852783
	pesos_i(4749) := b"0000000000000000_0000000000000000_0100101000010101_0111011100000000"; -- 0.28939002752304077
	pesos_i(4750) := b"0000000000000000_0000000000000000_0100110011111100_1111111110000000"; -- 0.3007354438304901
	pesos_i(4751) := b"0000000000000000_0000000000000000_0011110000101001_0101001000000000"; -- 0.23500549793243408
	pesos_i(4752) := b"0000000000000000_0000000000000000_0000000000001010_0000001010010011"; -- 0.00015274138422682881
	pesos_i(4753) := b"1111111111111111_1111111111111111_1101110011011101_1011011001000000"; -- -0.13724194467067719
	pesos_i(4754) := b"1111111111111111_1111111111111111_1011101100100100_1001000110000000"; -- -0.2689732611179352
	pesos_i(4755) := b"1111111111111111_1111111111111111_1111011000000000_0011110011010000"; -- -0.0390588752925396
	pesos_i(4756) := b"0000000000000000_0000000000000000_0011110100011000_1100100110000000"; -- 0.23865947127342224
	pesos_i(4757) := b"0000000000000000_0000000000000000_0010010100100011_0000011000000000"; -- 0.14506566524505615
	pesos_i(4758) := b"1111111111111111_1111111111111111_1110110000100110_0100001011100000"; -- -0.07754117995500565
	pesos_i(4759) := b"0000000000000000_0000000000000000_0001111001010101_0010011011000000"; -- 0.11848680675029755
	pesos_i(4760) := b"0000000000000000_0000000000000000_0100101011011000_1001111110000000"; -- 0.2923679053783417
	pesos_i(4761) := b"0000000000000000_0000000000000000_0011000010001011_0100010101000000"; -- 0.1896250993013382
	pesos_i(4762) := b"1111111111111111_1111111111111111_1111001100001101_0011001111100000"; -- -0.05057979375123978
	pesos_i(4763) := b"1111111111111111_1111111111111111_1100101011000011_0101011001000000"; -- -0.20795689523220062
	pesos_i(4764) := b"0000000000000000_0000000000000000_0001000101000111_1010111010100000"; -- 0.0675000324845314
	pesos_i(4765) := b"0000000000000000_0000000000000000_0010110110000111_1111010010000000"; -- 0.17785575985908508
	pesos_i(4766) := b"0000000000000000_0000000000000000_0011000011010111_1001111100000000"; -- 0.1907901167869568
	pesos_i(4767) := b"0000000000000000_0000000000000000_0010100110101100_0011101001000000"; -- 0.16278423368930817
	pesos_i(4768) := b"0000000000000000_0000000000000000_0000100110101111_0011101110110000"; -- 0.03783009573817253
	pesos_i(4769) := b"0000000000000000_0000000000000000_0010011100101011_1101000001000000"; -- 0.15301229059696198
	pesos_i(4770) := b"1111111111111111_1111111111111111_1110111011101010_1101011001000000"; -- -0.06672917306423187
	pesos_i(4771) := b"0000000000000000_0000000000000000_0000010101001101_0110110001010000"; -- 0.020712632685899734
	pesos_i(4772) := b"0000000000000000_0000000000000000_0001110001010111_0110100111000000"; -- 0.1107088178396225
	pesos_i(4773) := b"1111111111111111_1111111111111111_1100011010001101_1110100011000000"; -- -0.22439713776111603
	pesos_i(4774) := b"1111111111111111_1111111111111111_1101010011110101_1001000100000000"; -- -0.16812795400619507
	pesos_i(4775) := b"0000000000000000_0000000000000000_0011100100001011_1000111110000000"; -- 0.22283264994621277
	pesos_i(4776) := b"0000000000000000_0000000000000000_0101100100110101_1010000010000000"; -- 0.34847453236579895
	pesos_i(4777) := b"0000000000000000_0000000000000000_0000100011000001_0111001110010000"; -- 0.034201834350824356
	pesos_i(4778) := b"1111111111111111_1111111111111111_1011111000011000_0110110010000000"; -- -0.25743982195854187
	pesos_i(4779) := b"0000000000000000_0000000000000000_0000111101001010_0100110110110000"; -- 0.05972753092646599
	pesos_i(4780) := b"1111111111111111_1111111111111111_1111011000011100_0001001110000000"; -- -0.03863409161567688
	pesos_i(4781) := b"1111111111111111_1111111111111111_1100001000011010_0111101000000000"; -- -0.2417834997177124
	pesos_i(4782) := b"0000000000000000_0000000000000000_0100010010000100_1001101110000000"; -- 0.2676484286785126
	pesos_i(4783) := b"0000000000000000_0000000000000000_0010000110011000_0001110011000000"; -- 0.1312272995710373
	pesos_i(4784) := b"1111111111111111_1111111111111111_1001110111100011_1100011000000000"; -- -0.383243203163147
	pesos_i(4785) := b"1111111111111111_1111111111111111_1110110010000010_0010010100000000"; -- -0.07613915205001831
	pesos_i(4786) := b"1111111111111111_1111111111111111_1011100100011000_1000110100000000"; -- -0.27696913480758667
	pesos_i(4787) := b"0000000000000000_0000000000000000_0100011110011011_1111110110000000"; -- 0.27972397208213806
	pesos_i(4788) := b"0000000000000000_0000000000000000_0110111100010000_0101111110000000"; -- 0.43384358286857605
	pesos_i(4789) := b"1111111111111111_1111111111111111_1110111011001100_0101110100000000"; -- -0.06719416379928589
	pesos_i(4790) := b"1111111111111111_1111111111111111_0110011000110101_0010010000000000"; -- -0.6007516384124756
	pesos_i(4791) := b"0000000000000000_0000000000000000_0011101101101101_1001011000000000"; -- 0.2321408987045288
	pesos_i(4792) := b"1111111111111111_1111111111111111_1110110110000001_0010101011100000"; -- -0.07224781066179276
	pesos_i(4793) := b"0000000000000000_0000000000000000_0011101101011110_1101010111000000"; -- 0.23191581666469574
	pesos_i(4794) := b"0000000000000000_0000000000000000_0010010100100111_0110011100000000"; -- 0.14513248205184937
	pesos_i(4795) := b"1111111111111111_1111111111111111_1111010100100000_0001001001010000"; -- -0.04247937723994255
	pesos_i(4796) := b"1111111111111111_1111111111111111_1110100000011000_0100101100000000"; -- -0.09337931871414185
	pesos_i(4797) := b"1111111111111111_1111111111111111_1101010101011010_0110110101000000"; -- -0.1665889471769333
	pesos_i(4798) := b"0000000000000000_0000000000000000_0000101110001111_0000011001110000"; -- 0.04515114054083824
	pesos_i(4799) := b"0000000000000000_0000000000000000_0000100011001010_0011101011010000"; -- 0.03433578088879585
	pesos_i(4800) := b"0000000000000000_0000000000000000_0100110010111110_0111010100000000"; -- 0.2997811436653137
	pesos_i(4801) := b"1111111111111111_1111111111111111_1101011000010010_0000110100000000"; -- -0.16378706693649292
	pesos_i(4802) := b"1111111111111111_1111111111111111_1010010000010100_0001100110000000"; -- -0.3590683043003082
	pesos_i(4803) := b"1111111111111111_1111111111111111_1101100110101000_0110010000000000"; -- -0.14977431297302246
	pesos_i(4804) := b"0000000000000000_0000000000000000_0011011011010001_1101110000000000"; -- 0.21413969993591309
	pesos_i(4805) := b"1111111111111111_1111111111111111_1100110011111010_1001100001000000"; -- -0.19930122792720795
	pesos_i(4806) := b"1111111111111111_1111111111111111_1011100100001000_1100101110000000"; -- -0.2772095501422882
	pesos_i(4807) := b"0000000000000000_0000000000000000_0011100011111001_1110010000000000"; -- 0.2225630283355713
	pesos_i(4808) := b"0000000000000000_0000000000000000_0011000000111000_1111101011000000"; -- 0.18836943805217743
	pesos_i(4809) := b"1111111111111111_1111111111111111_1100011100111000_0001110001000000"; -- -0.2218000739812851
	pesos_i(4810) := b"1111111111111111_1111111111111111_1111001111011110_1110000010100000"; -- -0.04738041013479233
	pesos_i(4811) := b"0000000000000000_0000000000000000_0001000101010001_1000000001100000"; -- 0.06764986366033554
	pesos_i(4812) := b"1111111111111111_1111111111111111_1101011101101000_0001101001000000"; -- -0.15856777131557465
	pesos_i(4813) := b"0000000000000000_0000000000000000_1000100101101011_0111001000000000"; -- 0.5367957353591919
	pesos_i(4814) := b"1111111111111111_1111111111111111_1010011101001000_1011011100000000"; -- -0.3465467095375061
	pesos_i(4815) := b"1111111111111111_1111111111111111_1101100011011110_1011101011000000"; -- -0.1528514176607132
	pesos_i(4816) := b"0000000000000000_0000000000000000_0110001010101110_0100110010000000"; -- 0.3854720890522003
	pesos_i(4817) := b"0000000000000000_0000000000000000_0100111001111101_1001011000000000"; -- 0.3066037893295288
	pesos_i(4818) := b"0000000000000000_0000000000000000_0000001100001001_0101011100010000"; -- 0.011861268430948257
	pesos_i(4819) := b"0000000000000000_0000000000000000_0001111100001101_0000111000100000"; -- 0.12129295617341995
	pesos_i(4820) := b"0000000000000000_0000000000000000_0010110101101101_1110011001000000"; -- 0.17745818197727203
	pesos_i(4821) := b"0000000000000000_0000000000000000_0100010100111010_1001011000000000"; -- 0.2704252004623413
	pesos_i(4822) := b"0000000000000000_0000000000000000_0110011000011101_1001111100000000"; -- 0.3988894820213318
	pesos_i(4823) := b"0000000000000000_0000000000000000_0100100010011101_0110100010000000"; -- 0.28365185856819153
	pesos_i(4824) := b"0000000000000000_0000000000000000_0011111001111100_0011011111000000"; -- 0.24408291280269623
	pesos_i(4825) := b"0000000000000000_0000000000000000_0100110111100101_1111001010000000"; -- 0.30428996682167053
	pesos_i(4826) := b"0000000000000000_0000000000000000_0011011111111100_0110100001000000"; -- 0.21869517862796783
	pesos_i(4827) := b"0000000000000000_0000000000000000_0010011100011010_0000000101000000"; -- 0.15274055302143097
	pesos_i(4828) := b"0000000000000000_0000000000000000_0010111100111101_1101110111000000"; -- 0.18453775346279144
	pesos_i(4829) := b"0000000000000000_0000000000000000_0001101010001101_1100110110100000"; -- 0.10372624546289444
	pesos_i(4830) := b"0000000000000000_0000000000000000_0001011100011010_0101101100000000"; -- 0.09024590253829956
	pesos_i(4831) := b"0000000000000000_0000000000000000_0010001100111000_0100011100000000"; -- 0.13757747411727905
	pesos_i(4832) := b"1111111111111111_1111111111111111_1000110001110010_1111100110000000"; -- -0.45137062668800354
	pesos_i(4833) := b"0000000000000000_0000000000000000_0000011001001010_0000110000110000"; -- 0.0245673768222332
	pesos_i(4834) := b"0000000000000000_0000000000000000_0001001000001111_1000111011100000"; -- 0.07054989784955978
	pesos_i(4835) := b"0000000000000000_0000000000000000_0010110000001110_0110111111000000"; -- 0.17209528386592865
	pesos_i(4836) := b"0000000000000000_0000000000000000_0001110100100000_1010111001000000"; -- 0.11377991735935211
	pesos_i(4837) := b"1111111111111111_1111111111111111_1100011100101011_1111101110000000"; -- -0.2219851315021515
	pesos_i(4838) := b"1111111111111111_1111111111111111_1011101101000000_1111010110000000"; -- -0.26854005455970764
	pesos_i(4839) := b"1111111111111111_1111111111111111_1010100100000110_1011011000000000"; -- -0.3397413492202759
	pesos_i(4840) := b"0000000000000000_0000000000000000_0001110001010111_1010100000000000"; -- 0.11071252822875977
	pesos_i(4841) := b"0000000000000000_0000000000000000_0100011111100001_0000101000000000"; -- 0.28077757358551025
	pesos_i(4842) := b"0000000000000000_0000000000000000_0011100100111011_0001100111000000"; -- 0.22355805337429047
	pesos_i(4843) := b"0000000000000000_0000000000000000_0001111110101001_0101101011000000"; -- 0.12367789447307587
	pesos_i(4844) := b"0000000000000000_0000000000000000_0011011100001011_0110010111000000"; -- 0.2150176614522934
	pesos_i(4845) := b"0000000000000000_0000000000000000_0111001001001100_1111110100000000"; -- 0.4464872479438782
	pesos_i(4846) := b"1111111111111111_1111111111111111_1111110000100001_1110011000110000"; -- -0.015107739716768265
	pesos_i(4847) := b"1111111111111111_1111111111111111_1101110000111010_0011101101000000"; -- -0.13973645865917206
	pesos_i(4848) := b"1111111111111111_1111111111111111_1100100101001111_0110000110000000"; -- -0.2136324942111969
	pesos_i(4849) := b"1111111111111111_1111111111111111_1110111010010001_1101011111000000"; -- -0.06808711588382721
	pesos_i(4850) := b"0000000000000000_0000000000000000_0101101010110111_1011111000000000"; -- 0.3543661832809448
	pesos_i(4851) := b"0000000000000000_0000000000000000_1000110110001101_1101010100000000"; -- 0.5529454350471497
	pesos_i(4852) := b"1111111111111111_1111111111111111_1110110000010111_1111100000100000"; -- -0.0777592584490776
	pesos_i(4853) := b"0000000000000000_0000000000000000_0011000000001110_0111010010000000"; -- 0.18772056698799133
	pesos_i(4854) := b"0000000000000000_0000000000000000_0100111010010101_0100000100000000"; -- 0.3069649338722229
	pesos_i(4855) := b"0000000000000000_0000000000000000_0000011100100000_0010101101101000"; -- 0.027834618464112282
	pesos_i(4856) := b"0000000000000000_0000000000000000_0010011111011110_1001011111000000"; -- 0.15574024617671967
	pesos_i(4857) := b"0000000000000000_0000000000000000_0011010100110100_1100111011000000"; -- 0.2078370302915573
	pesos_i(4858) := b"1111111111111111_1111111111111111_1111000000001001_1110110100100000"; -- -0.062348537147045135
	pesos_i(4859) := b"0000000000000000_0000000000000000_0001110010101010_0001110000100000"; -- 0.11197067052125931
	pesos_i(4860) := b"1111111111111111_1111111111111111_1010101010000000_1101101110000000"; -- -0.3339712917804718
	pesos_i(4861) := b"0000000000000000_0000000000000000_0011100101111110_1001010110000000"; -- 0.22458776831626892
	pesos_i(4862) := b"1111111111111111_1111111111111111_1010101110000011_0110100010000000"; -- -0.33002611994743347
	pesos_i(4863) := b"1111111111111111_1111111111111111_1111100001101110_0100000101000000"; -- -0.029567644000053406
	pesos_i(4864) := b"0000000000000000_0000000000000000_0010011101000011_1000001100000000"; -- 0.15337389707565308
	pesos_i(4865) := b"0000000000000000_0000000000000000_0010110001110101_0011000010000000"; -- 0.1736631691455841
	pesos_i(4866) := b"1111111111111111_1111111111111111_1101001010011110_1110111100000000"; -- -0.17726236581802368
	pesos_i(4867) := b"0000000000000000_0000000000000000_0010010011000101_1001111011000000"; -- 0.1436404436826706
	pesos_i(4868) := b"1111111111111111_1111111111111111_1111100010010000_1101001000010000"; -- -0.02904021367430687
	pesos_i(4869) := b"1111111111111111_1111111111111111_0111011011110011_0100010000000000"; -- -0.5353505611419678
	pesos_i(4870) := b"1111111111111111_1111111111111111_1111011110110101_0110001000110000"; -- -0.032388556748628616
	pesos_i(4871) := b"0000000000000000_0000000000000000_0011010001111101_1101010111000000"; -- 0.20504508912563324
	pesos_i(4872) := b"1111111111111111_1111111111111111_1110100110100110_1111101111100000"; -- -0.0872957780957222
	pesos_i(4873) := b"1111111111111111_1111111111111111_1111001111011111_0111001000100000"; -- -0.04737173765897751
	pesos_i(4874) := b"1111111111111111_1111111111111111_1111000110001000_1000110011110000"; -- -0.05651015415787697
	pesos_i(4875) := b"0000000000000000_0000000000000000_0000101001100100_1111111001000000"; -- 0.04060353338718414
	pesos_i(4876) := b"0000000000000000_0000000000000000_0001010100001001_1010101101000000"; -- 0.08217878639698029
	pesos_i(4877) := b"0000000000000000_0000000000000000_0000100010100101_0101101011010000"; -- 0.033773113042116165
	pesos_i(4878) := b"0000000000000000_0000000000000000_0100001000101011_1100001000000000"; -- 0.2584801912307739
	pesos_i(4879) := b"0000000000000000_0000000000000000_0010001100111000_1000100101000000"; -- 0.13758142292499542
	pesos_i(4880) := b"0000000000000000_0000000000000000_0000001000001010_0110101010001100"; -- 0.007971438579261303
	pesos_i(4881) := b"0000000000000000_0000000000000000_0001010100101010_1011010100000000"; -- 0.08268290758132935
	pesos_i(4882) := b"1111111111111111_1111111111111111_1110000010001001_0100011110000000"; -- -0.12290528416633606
	pesos_i(4883) := b"1111111111111111_1111111111111111_1111111110011110_1100000001111010"; -- -0.001483888947404921
	pesos_i(4884) := b"0000000000000000_0000000000000000_0011011000011101_1111001111000000"; -- 0.2113945335149765
	pesos_i(4885) := b"1111111111111111_1111111111111111_1110010100100110_1100111000100000"; -- -0.10487663000822067
	pesos_i(4886) := b"0000000000000000_0000000000000000_0011000000101110_0101111100000000"; -- 0.18820756673812866
	pesos_i(4887) := b"1111111111111111_1111111111111111_1111101000110111_1101011011110000"; -- -0.02258545532822609
	pesos_i(4888) := b"0000000000000000_0000000000000000_0011110000111011_0111111001000000"; -- 0.2352827936410904
	pesos_i(4889) := b"0000000000000000_0000000000000000_0001011100111010_1011110101000000"; -- 0.09074003994464874
	pesos_i(4890) := b"0000000000000000_0000000000000000_0000000000101100_0110011000111001"; -- 0.0006774796056561172
	pesos_i(4891) := b"1111111111111111_1111111111111111_1111110110011111_0111010111000100"; -- -0.009285583160817623
	pesos_i(4892) := b"0000000000000000_0000000000000000_0001100000111011_0001000010100000"; -- 0.09465125948190689
	pesos_i(4893) := b"0000000000000000_0000000000000000_0100100101101110_0110011000000000"; -- 0.2868407964706421
	pesos_i(4894) := b"0000000000000000_0000000000000000_0100001001111001_1110010000000000"; -- 0.2596724033355713
	pesos_i(4895) := b"1111111111111111_1111111111111111_1110100101101110_1111110010000000"; -- -0.08815023303031921
	pesos_i(4896) := b"0000000000000000_0000000000000000_0010011100001101_0001100010000000"; -- 0.1525435745716095
	pesos_i(4897) := b"0000000000000000_0000000000000000_0011000010101110_1101111111000000"; -- 0.1901683658361435
	pesos_i(4898) := b"0000000000000000_0000000000000000_0011100000111001_0110110101000000"; -- 0.2196262627840042
	pesos_i(4899) := b"0000000000000000_0000000000000000_0010000101100000_1101001010000000"; -- 0.13038364052772522
	pesos_i(4900) := b"1111111111111111_1111111111111111_1011100100000001_0100111000000000"; -- -0.277323842048645
	pesos_i(4901) := b"0000000000000000_0000000000000000_0000001011111100_0010110011001100"; -- 0.011660384945571423
	pesos_i(4902) := b"1111111111111111_1111111111111111_1111000011011101_1010100110000000"; -- -0.05911770462989807
	pesos_i(4903) := b"0000000000000000_0000000000000000_0011010111101011_0110110110000000"; -- 0.2106235921382904
	pesos_i(4904) := b"1111111111111111_1111111111111111_1110101010101010_0111000011100000"; -- -0.08333677798509598
	pesos_i(4905) := b"1111111111111111_1111111111111111_1111000001000010_1010011011110000"; -- -0.06148296967148781
	pesos_i(4906) := b"0000000000000000_0000000000000000_0010100001000000_0000110101000000"; -- 0.15722735226154327
	pesos_i(4907) := b"1111111111111111_1111111111111111_1100101100010111_0000110101000000"; -- -0.20667950809001923
	pesos_i(4908) := b"0000000000000000_0000000000000000_0011010101001100_1011001101000000"; -- 0.208201602101326
	pesos_i(4909) := b"1111111111111111_1111111111111111_1011010010010010_1010100000000000"; -- -0.29463720321655273
	pesos_i(4910) := b"1111111111111111_1111111111111111_1110101001010001_0000011100100000"; -- -0.08470111340284348
	pesos_i(4911) := b"0000000000000000_0000000000000000_0000111010000110_0000010001100000"; -- 0.05673243850469589
	pesos_i(4912) := b"1111111111111111_1111111111111111_1100111011110111_0001111000000000"; -- -0.19154179096221924
	pesos_i(4913) := b"0000000000000000_0000000000000000_0011111100010000_0000111100000000"; -- 0.24633878469467163
	pesos_i(4914) := b"1111111111111111_1111111111111111_1001100001101111_0010100000000000"; -- -0.4045538902282715
	pesos_i(4915) := b"0000000000000000_0000000000000000_0001001000110111_1111010001000000"; -- 0.07116629183292389
	pesos_i(4916) := b"0000000000000000_0000000000000000_0010110101011011_1111010011000000"; -- 0.17718438804149628
	pesos_i(4917) := b"1111111111111111_1111111111111111_1111101110111001_1110100100001000"; -- -0.016694484278559685
	pesos_i(4918) := b"1111111111111111_1111111111111111_1001010101001100_0111010000000000"; -- -0.41680216789245605
	pesos_i(4919) := b"0000000000000000_0000000000000000_0000111110011110_0111101100000000"; -- 0.06101197004318237
	pesos_i(4920) := b"0000000000000000_0000000000000000_0001001010010111_0000101000100000"; -- 0.07261718064546585
	pesos_i(4921) := b"0000000000000000_0000000000000000_0010100110110111_0001101101000000"; -- 0.16295023262500763
	pesos_i(4922) := b"0000000000000000_0000000000000000_0000110000010000_1101011010010000"; -- 0.04713192954659462
	pesos_i(4923) := b"0000000000000000_0000000000000000_0001011001110110_1101110110100000"; -- 0.08775124698877335
	pesos_i(4924) := b"1111111111111111_1111111111111111_1110101010100111_0010011110000000"; -- -0.08338692784309387
	pesos_i(4925) := b"0000000000000000_0000000000000000_0001101101001101_1000000000100000"; -- 0.10665131360292435
	pesos_i(4926) := b"0000000000000000_0000000000000000_0000001101001011_0100100011100000"; -- 0.012867502868175507
	pesos_i(4927) := b"0000000000000000_0000000000000000_0010001010111100_1111000101000000"; -- 0.13569553196430206
	pesos_i(4928) := b"1111111111111111_1111111111111111_1100110010010111_1000001000000000"; -- -0.2008131742477417
	pesos_i(4929) := b"1111111111111111_1111111111111111_1011101001011101_1110100010000000"; -- -0.2720045745372772
	pesos_i(4930) := b"1111111111111111_1111111111111111_1100111000011111_0101000011000000"; -- -0.1948346644639969
	pesos_i(4931) := b"1111111111111111_1111111111111111_1101100101000110_1110010000000000"; -- -0.1512620449066162
	pesos_i(4932) := b"0000000000000000_0000000000000000_0001000000011000_0001100101100000"; -- 0.06286772340536118
	pesos_i(4933) := b"0000000000000000_0000000000000000_0000010101101100_1101111101000000"; -- 0.021192505955696106
	pesos_i(4934) := b"1111111111111111_1111111111111111_1001100100100110_1101101110000000"; -- -0.4017508327960968
	pesos_i(4935) := b"1111111111111111_1111111111111111_1011111111000010_1101001000000000"; -- -0.25093352794647217
	pesos_i(4936) := b"0000000000000000_0000000000000000_0000010111001101_0101000111011000"; -- 0.022664180025458336
	pesos_i(4937) := b"1111111111111111_1111111111111111_1101011011000000_1001011000000000"; -- -0.1611238718032837
	pesos_i(4938) := b"1111111111111111_1111111111111111_1111111110100100_1011011010001110"; -- -0.0013929273700341582
	pesos_i(4939) := b"0000000000000000_0000000000000000_0010110110010110_1011110000000000"; -- 0.17808127403259277
	pesos_i(4940) := b"1111111111111111_1111111111111111_1010011100010011_1100100110000000"; -- -0.34735432267189026
	pesos_i(4941) := b"1111111111111111_1111111111111111_1110111110101100_0110000110100000"; -- -0.0637759193778038
	pesos_i(4942) := b"1111111111111111_1111111111111111_1100011000001101_1001110000000000"; -- -0.22635483741760254
	pesos_i(4943) := b"1111111111111111_1111111111111111_1111100110010100_0110011100100000"; -- -0.025079302489757538
	pesos_i(4944) := b"0000000000000000_0000000000000000_0010000110001001_1010011010000000"; -- 0.1310066282749176
	pesos_i(4945) := b"0000000000000000_0000000000000000_0100100111100011_1010010010000000"; -- 0.28862980008125305
	pesos_i(4946) := b"0000000000000000_0000000000000000_0001011101000111_0011101010000000"; -- 0.09093061089515686
	pesos_i(4947) := b"0000000000000000_0000000000000000_0001111000000000_0110001110100000"; -- 0.11719343811273575
	pesos_i(4948) := b"0000000000000000_0000000000000000_0001101101110100_1110000100100000"; -- 0.10725218802690506
	pesos_i(4949) := b"1111111111111111_1111111111111111_1110100000000000_1011001000100000"; -- -0.09373938292264938
	pesos_i(4950) := b"0000000000000000_0000000000000000_0011000011000000_1000110110000000"; -- 0.19043812155723572
	pesos_i(4951) := b"1111111111111111_1111111111111111_1110101001111101_0000111101000000"; -- -0.08402924239635468
	pesos_i(4952) := b"0000000000000000_0000000000000000_0010011100001000_0101000101000000"; -- 0.152470663189888
	pesos_i(4953) := b"0000000000000000_0000000000000000_0000001011100101_0111101001010000"; -- 0.01131405308842659
	pesos_i(4954) := b"1111111111111111_1111111111111111_1101101101100000_1011010110000000"; -- -0.14305558800697327
	pesos_i(4955) := b"1111111111111111_1111111111111111_1111010001111101_1110011000000000"; -- -0.04495394229888916
	pesos_i(4956) := b"0000000000000000_0000000000000000_0100000100110111_0100000110000000"; -- 0.2547493875026703
	pesos_i(4957) := b"1111111111111111_1111111111111111_1100010111101101_1110111111000000"; -- -0.2268381267786026
	pesos_i(4958) := b"0000000000000000_0000000000000000_0010100110001111_0000101110000000"; -- 0.16233894228935242
	pesos_i(4959) := b"0000000000000000_0000000000000000_0000101100011101_0100010110110000"; -- 0.043415408581495285
	pesos_i(4960) := b"1111111111111111_1111111111111111_0111111000000011_1111001000000000"; -- -0.5077522993087769
	pesos_i(4961) := b"1111111111111111_1111111111111111_1101101110101000_1100110001000000"; -- -0.14195559918880463
	pesos_i(4962) := b"1111111111111111_1111111111111111_1100011011110100_0101000000000000"; -- -0.22283458709716797
	pesos_i(4963) := b"1111111111111111_1111111111111111_1111011100110101_1001110100000000"; -- -0.034338176250457764
	pesos_i(4964) := b"1111111111111111_1111111111111111_1110011110011100_1001101010100000"; -- -0.0952666625380516
	pesos_i(4965) := b"0000000000000000_0000000000000000_0001110000110001_0010101111000000"; -- 0.11012528836727142
	pesos_i(4966) := b"0000000000000000_0000000000000000_0000101110100100_1000111000000000"; -- 0.045479655265808105
	pesos_i(4967) := b"1111111111111111_1111111111111111_0110100001100000_1000011100000000"; -- -0.5922771096229553
	pesos_i(4968) := b"1111111111111111_1111111111111111_1110001100101111_0110101100000000"; -- -0.11255770921707153
	pesos_i(4969) := b"1111111111111111_1111111111111111_1110100011010110_1000110100100000"; -- -0.09047620743513107
	pesos_i(4970) := b"0000000000000000_0000000000000000_0000101000011010_0101101011010000"; -- 0.039464641362428665
	pesos_i(4971) := b"0000000000000000_0000000000000000_0000110000011101_0001011010110000"; -- 0.04731885716319084
	pesos_i(4972) := b"0000000000000000_0000000000000000_0001011111111001_0110011001100000"; -- 0.09364929050207138
	pesos_i(4973) := b"1111111111111111_1111111111111111_1100110100010110_1011100110000000"; -- -0.19887199997901917
	pesos_i(4974) := b"1111111111111111_1111111111111111_1101001111100111_0100101100000000"; -- -0.17225199937820435
	pesos_i(4975) := b"1111111111111111_1111111111111111_1011101111101101_1101011010000000"; -- -0.2659021317958832
	pesos_i(4976) := b"1111111111111111_1111111111111111_1111101100000000_1100001101111000"; -- -0.01951959915459156
	pesos_i(4977) := b"0000000000000000_0000000000000000_0010000001100011_1111100100000000"; -- 0.12652546167373657
	pesos_i(4978) := b"0000000000000000_0000000000000000_0110011010000110_0111001110000000"; -- 0.40048906207084656
	pesos_i(4979) := b"0000000000000000_0000000000000000_0000100100000010_0001010111100000"; -- 0.03518807142972946
	pesos_i(4980) := b"0000000000000000_0000000000000000_0001011000101011_1101101101100000"; -- 0.0866067036986351
	pesos_i(4981) := b"0000000000000000_0000000000000000_0001011100011111_1101100101000000"; -- 0.09032972157001495
	pesos_i(4982) := b"0000000000000000_0000000000000000_0010110011110110_1100011011000000"; -- 0.1756405085325241
	pesos_i(4983) := b"0000000000000000_0000000000000000_0001010011110100_0111011100100000"; -- 0.08185524493455887
	pesos_i(4984) := b"0000000000000000_0000000000000000_0001101110011110_1001000000100000"; -- 0.10788822919130325
	pesos_i(4985) := b"0000000000000000_0000000000000000_0000100110010101_0010010010010000"; -- 0.0374319888651371
	pesos_i(4986) := b"1111111111111111_1111111111111111_1110010101101101_0100101000000000"; -- -0.10380113124847412
	pesos_i(4987) := b"1111111111111111_1111111111111111_1101110100000011_0110111001000000"; -- -0.136666402220726
	pesos_i(4988) := b"0000000000000000_0000000000000000_0001010110101011_0110001001100000"; -- 0.08464636653661728
	pesos_i(4989) := b"1111111111111111_1111111111111111_1110111000011100_1001111011000000"; -- -0.0698757916688919
	pesos_i(4990) := b"1111111111111111_1111111111111111_1011010011100110_0010111100000000"; -- -0.29336267709732056
	pesos_i(4991) := b"1111111111111111_1111111111111111_1001010110111111_1101010010000000"; -- -0.41504165530204773
	pesos_i(4992) := b"0000000000000000_0000000000000000_0000100110001100_0010001100000000"; -- 0.03729456663131714
	pesos_i(4993) := b"0000000000000000_0000000000000000_0011110110001011_1110011110000000"; -- 0.240416020154953
	pesos_i(4994) := b"1111111111111111_1111111111111111_1111101101010110_0011010101101000"; -- -0.018215810880064964
	pesos_i(4995) := b"0000000000000000_0000000000000000_0001000011101101_1000011111000000"; -- 0.06612442433834076
	pesos_i(4996) := b"0000000000000000_0000000000000000_0000101000011010_1100000011110000"; -- 0.03947072848677635
	pesos_i(4997) := b"0000000000000000_0000000000000000_0001011100000010_1010110110000000"; -- 0.08988460898399353
	pesos_i(4998) := b"0000000000000000_0000000000000000_0100010001011111_1001110110000000"; -- 0.2670839726924896
	pesos_i(4999) := b"0000000000000000_0000000000000000_0000110110000101_0111000100110000"; -- 0.052817415446043015
	pesos_i(5000) := b"0000000000000000_0000000000000000_0000110101010011_1101110110000000"; -- 0.05206093192100525
	pesos_i(5001) := b"0000000000000000_0000000000000000_0100100001110001_0111000100000000"; -- 0.2829809784889221
	pesos_i(5002) := b"1111111111111111_1111111111111111_1110101011001100_1110001110000000"; -- -0.0828111469745636
	pesos_i(5003) := b"1111111111111111_1111111111111111_1111101011111110_1101110010000000"; -- -0.019548624753952026
	pesos_i(5004) := b"1111111111111111_1111111111111111_1110110000110011_1110110001100000"; -- -0.07733271270990372
	pesos_i(5005) := b"0000000000000000_0000000000000000_0010101001010010_0111111001000000"; -- 0.1653212457895279
	pesos_i(5006) := b"0000000000000000_0000000000000000_0001001001100110_1000000000100000"; -- 0.07187653332948685
	pesos_i(5007) := b"1111111111111111_1111111111111111_1110111000011001_0110000110100000"; -- -0.0699252113699913
	pesos_i(5008) := b"1111111111111111_1111111111111111_1110011110011111_1111101101100000"; -- -0.09521511942148209
	pesos_i(5009) := b"0000000000000000_0000000000000000_0100101011011001_1101111010000000"; -- 0.292386919260025
	pesos_i(5010) := b"1111111111111111_1111111111111111_1110000001101111_1101110000000000"; -- -0.12329316139221191
	pesos_i(5011) := b"0000000000000000_0000000000000000_0011011110110101_1111110011000000"; -- 0.21762065589427948
	pesos_i(5012) := b"0000000000000000_0000000000000000_0001110010111111_1110000010100000"; -- 0.11230281740427017
	pesos_i(5013) := b"0000000000000000_0000000000000000_0001000011100010_0000010001000000"; -- 0.0659487396478653
	pesos_i(5014) := b"0000000000000000_0000000000000000_0011111010010111_0110010001000000"; -- 0.24449755251407623
	pesos_i(5015) := b"1111111111111111_1111111111111111_1101000111110101_0001101000000000"; -- -0.17985379695892334
	pesos_i(5016) := b"0000000000000000_0000000000000000_0011000100000110_0011011110000000"; -- 0.19150111079216003
	pesos_i(5017) := b"1111111111111111_1111111111111111_1100011011111001_1110001001000000"; -- -0.22274957597255707
	pesos_i(5018) := b"1111111111111111_1111111111111111_1111111011010100_1111110100101010"; -- -0.004562546964734793
	pesos_i(5019) := b"0000000000000000_0000000000000000_0000111010001010_1011110111010000"; -- 0.05680452659726143
	pesos_i(5020) := b"1111111111111111_1111111111111111_1111110111100101_1111001101000100"; -- -0.008209987543523312
	pesos_i(5021) := b"0000000000000000_0000000000000000_0011111101000010_0000111011000000"; -- 0.24710170924663544
	pesos_i(5022) := b"0000000000000000_0000000000000000_0011001000001100_0111000111000000"; -- 0.1955023854970932
	pesos_i(5023) := b"0000000000000000_0000000000000000_0010011001011101_1011001011000000"; -- 0.1498672217130661
	pesos_i(5024) := b"0000000000000000_0000000000000000_0001011111001010_0011010001000000"; -- 0.09292913973331451
	pesos_i(5025) := b"0000000000000000_0000000000000000_0001110110111010_1110000111000000"; -- 0.11613284051418304
	pesos_i(5026) := b"0000000000000000_0000000000000000_0000100011110001_1101000000100000"; -- 0.03493977338075638
	pesos_i(5027) := b"0000000000000000_0000000000000000_0000001100000011_0001001010111100"; -- 0.011765643022954464
	pesos_i(5028) := b"1111111111111111_1111111111111111_1011000001101000_1111001100000000"; -- -0.3108986020088196
	pesos_i(5029) := b"0000000000000000_0000000000000000_0001101100101101_0101111010000000"; -- 0.10616102814674377
	pesos_i(5030) := b"1111111111111111_1111111111111111_1101110000100001_1100011111000000"; -- -0.14010955393314362
	pesos_i(5031) := b"1111111111111111_1111111111111111_1101110010001111_1101000111000000"; -- -0.13843049108982086
	pesos_i(5032) := b"1111111111111111_1111111111111111_1100000111011001_1000101101000000"; -- -0.24277429282665253
	pesos_i(5033) := b"1111111111111111_1111111111111111_1110100111010001_0010000000000000"; -- -0.08665275573730469
	pesos_i(5034) := b"0000000000000000_0000000000000000_0000011000101111_0100011000110000"; -- 0.024158846586942673
	pesos_i(5035) := b"1111111111111111_1111111111111111_1011111110000001_0101011010000000"; -- -0.25193271040916443
	pesos_i(5036) := b"0000000000000000_0000000000000000_0010111110100010_0010011011000000"; -- 0.18606798350811005
	pesos_i(5037) := b"0000000000000000_0000000000000000_0000100100100100_0011001010100000"; -- 0.035708583891391754
	pesos_i(5038) := b"1111111111111111_1111111111111111_1110011101010011_1100101110000000"; -- -0.09637764096260071
	pesos_i(5039) := b"0000000000000000_0000000000000000_0010001101011101_1110110001000000"; -- 0.13815189898014069
	pesos_i(5040) := b"1111111111111111_1111111111111111_1011010110011010_1001101000000000"; -- -0.2906097173690796
	pesos_i(5041) := b"0000000000000000_0000000000000000_0011010010011000_1000001110000000"; -- 0.20545217394828796
	pesos_i(5042) := b"1111111111111111_1111111111111111_1101110101000010_1100000110000000"; -- -0.13570013642311096
	pesos_i(5043) := b"1111111111111111_1111111111111111_1111001010110110_1110000100000000"; -- -0.05189698934555054
	pesos_i(5044) := b"0000000000000000_0000000000000000_0000001011010101_0111000100011100"; -- 0.011069363914430141
	pesos_i(5045) := b"1111111111111111_1111111111111111_1110001100100010_0001101010100000"; -- -0.11276086419820786
	pesos_i(5046) := b"1111111111111111_1111111111111111_1100001100000101_0000010000000000"; -- -0.2382047176361084
	pesos_i(5047) := b"0000000000000000_0000000000000000_0011110111100110_0000101011000000"; -- 0.24179141223430634
	pesos_i(5048) := b"1111111111111111_1111111111111111_1011101101001000_0101110010000000"; -- -0.2684271037578583
	pesos_i(5049) := b"1111111111111111_1111111111111111_1110011000101110_0000000011000000"; -- -0.10086055099964142
	pesos_i(5050) := b"1111111111111111_1111111111111111_1100010000011000_0101111111000000"; -- -0.23400308191776276
	pesos_i(5051) := b"0000000000000000_0000000000000000_0001010101111010_1011000011100000"; -- 0.08390336483716965
	pesos_i(5052) := b"1111111111111111_1111111111111111_1100111111000100_0000100011000000"; -- -0.18841500580310822
	pesos_i(5053) := b"1111111111111111_1111111111111111_1110101010100111_0000111001000000"; -- -0.08338843286037445
	pesos_i(5054) := b"1111111111111111_1111111111111111_1111111011101100_0110100010010000"; -- -0.004205193370580673
	pesos_i(5055) := b"0000000000000000_0000000000000000_0000000110011000_0110011111010100"; -- 0.00623177457600832
	pesos_i(5056) := b"1111111111111111_1111111111111111_1111001110000001_0010000110100000"; -- -0.04881086200475693
	pesos_i(5057) := b"1111111111111111_1111111111111111_1001000001101000_1101100000000000"; -- -0.4359002113342285
	pesos_i(5058) := b"0000000000000000_0000000000000000_0001001010111101_1001001001100000"; -- 0.0732051357626915
	pesos_i(5059) := b"1111111111111111_1111111111111111_1110001101010010_0111101110100000"; -- -0.11202266067266464
	pesos_i(5060) := b"1111111111111111_1111111111111111_1100010101001010_1110010000000000"; -- -0.2293260097503662
	pesos_i(5061) := b"0000000000000000_0000000000000000_0100001010111001_0000000100000000"; -- 0.2606354355812073
	pesos_i(5062) := b"1111111111111111_1111111111111111_1110000100111101_0110000100100000"; -- -0.12015717476606369
	pesos_i(5063) := b"1111111111111111_1111111111111111_1101110110111010_1010000000000000"; -- -0.13387107849121094
	pesos_i(5064) := b"0000000000000000_0000000000000000_0000010001110001_1111111000000000"; -- 0.01736438274383545
	pesos_i(5065) := b"1111111111111111_1111111111111111_1100001101010111_0010100110000000"; -- -0.23695126175880432
	pesos_i(5066) := b"1111111111111111_1111111111111111_1010111100001101_1000001010000000"; -- -0.3162001073360443
	pesos_i(5067) := b"1111111111111111_1111111111111111_1110100001010001_0101000010000000"; -- -0.09250923991203308
	pesos_i(5068) := b"1111111111111111_1111111111111111_1100011001110100_0001111101000000"; -- -0.22479061782360077
	pesos_i(5069) := b"1111111111111111_1111111111111111_1111011011010101_0010111001100000"; -- -0.03580961376428604
	pesos_i(5070) := b"1111111111111111_1111111111111111_1111010111001101_0100001110100000"; -- -0.039836667478084564
	pesos_i(5071) := b"1111111111111111_1111111111111111_1101010000110001_0011111101000000"; -- -0.17112354934215546
	pesos_i(5072) := b"1111111111111111_1111111111111111_1101011110000111_0011111110000000"; -- -0.15809252858161926
	pesos_i(5073) := b"1111111111111111_1111111111111111_1101110011010000_1010011010000000"; -- -0.1374412477016449
	pesos_i(5074) := b"0000000000000000_0000000000000000_0010010110011101_1000110000000000"; -- 0.14693522453308105
	pesos_i(5075) := b"0000000000000000_0000000000000000_0100011000111111_0101100000000000"; -- 0.27440404891967773
	pesos_i(5076) := b"0000000000000000_0000000000000000_0001000111101111_1111001101000000"; -- 0.07006759941577911
	pesos_i(5077) := b"1111111111111111_1111111111111111_1111000010001010_0111010011110000"; -- -0.06038731709122658
	pesos_i(5078) := b"0000000000000000_0000000000000000_0001011101100010_0010101011000000"; -- 0.09134165942668915
	pesos_i(5079) := b"1111111111111111_1111111111111111_1111011011110001_1111111101100000"; -- -0.035369910299777985
	pesos_i(5080) := b"0000000000000000_0000000000000000_0001101101110110_1001111000100000"; -- 0.10727871209383011
	pesos_i(5081) := b"0000000000000000_0000000000000000_0000110001001000_1000010000010000"; -- 0.04798150435090065
	pesos_i(5082) := b"1111111111111111_1111111111111111_1110100010000010_0110110010100000"; -- -0.09175988286733627
	pesos_i(5083) := b"0000000000000000_0000000000000000_0000110000111001_0010101011000000"; -- 0.04774729907512665
	pesos_i(5084) := b"0000000000000000_0000000000000000_0001111010000101_1010111110000000"; -- 0.11922737956047058
	pesos_i(5085) := b"1111111111111111_1111111111111111_1010111110100101_1111000000000000"; -- -0.3138742446899414
	pesos_i(5086) := b"1111111111111111_1111111111111111_1100101111111110_0000000001000000"; -- -0.2031555026769638
	pesos_i(5087) := b"0000000000000000_0000000000000000_0010101110101001_1100101001000000"; -- 0.17055954039096832
	pesos_i(5088) := b"1111111111111111_1111111111111111_1011011001111110_1111010110000000"; -- -0.28712525963783264
	pesos_i(5089) := b"0000000000000000_0000000000000000_0010000101000010_0011111111000000"; -- 0.12991712987422943
	pesos_i(5090) := b"1111111111111111_1111111111111111_1111010101000111_1000111000010000"; -- -0.041876908391714096
	pesos_i(5091) := b"1111111111111111_1111111111111111_1101101101111111_1000001110000000"; -- -0.14258554577827454
	pesos_i(5092) := b"1111111111111111_1111111111111111_1111111011100010_0101011001100110"; -- -0.004358863923698664
	pesos_i(5093) := b"1111111111111111_1111111111111111_1010100011110100_0111000110000000"; -- -0.340020090341568
	pesos_i(5094) := b"0000000000000000_0000000000000000_0010011011000101_1011000110000000"; -- 0.15145406126976013
	pesos_i(5095) := b"1111111111111111_1111111111111111_1001111010111010_1100111110000000"; -- -0.3799619972705841
	pesos_i(5096) := b"1111111111111111_1111111111111111_1100000111000001_1101011101000000"; -- -0.2431359738111496
	pesos_i(5097) := b"1111111111111111_1111111111111111_0111010010000001_1110110100000000"; -- -0.5448924899101257
	pesos_i(5098) := b"0000000000000000_0000000000000000_0000100100100001_0001110001000000"; -- 0.035661473870277405
	pesos_i(5099) := b"0000000000000000_0000000000000000_0011000010010001_1101110010000000"; -- 0.18972566723823547
	pesos_i(5100) := b"0000000000000000_0000000000000000_0011001110111101_1010000011000000"; -- 0.20211224257946014
	pesos_i(5101) := b"1111111111111111_1111111111111111_1001011001001110_1101100110000000"; -- -0.41285935044288635
	pesos_i(5102) := b"0000000000000000_0000000000000000_0000011111100001_1011011001110000"; -- 0.03078785166144371
	pesos_i(5103) := b"0000000000000000_0000000000000000_0010110100011111_0011110101000000"; -- 0.17625792324543
	pesos_i(5104) := b"0000000000000000_0000000000000000_0100100111101101_1101000010000000"; -- 0.28878501057624817
	pesos_i(5105) := b"0000000000000000_0000000000000000_0010011001101001_1101010011000000"; -- 0.15005235373973846
	pesos_i(5106) := b"0000000000000000_0000000000000000_0010110011101000_0111111110000000"; -- 0.17542263865470886
	pesos_i(5107) := b"0000000000000000_0000000000000000_0001001001011100_0110101110000000"; -- 0.07172271609306335
	pesos_i(5108) := b"1111111111111111_1111111111111111_1110011010000010_1000010000000000"; -- -0.09957098960876465
	pesos_i(5109) := b"1111111111111111_1111111111111111_1010100111110100_0001111010000000"; -- -0.33611878752708435
	pesos_i(5110) := b"0000000000000000_0000000000000000_0001110111011011_1110100110000000"; -- 0.11663684248924255
	pesos_i(5111) := b"0000000000000000_0000000000000000_0000001000001111_0110001100010100"; -- 0.008047287352383137
	pesos_i(5112) := b"0000000000000000_0000000000000000_0100001000011101_1000001000000000"; -- 0.2582627534866333
	pesos_i(5113) := b"1111111111111111_1111111111111111_1111001101110011_0110101100100000"; -- -0.049020104110240936
	pesos_i(5114) := b"0000000000000000_0000000000000000_0000101110101111_1111011011100000"; -- 0.045653752982616425
	pesos_i(5115) := b"1111111111111111_1111111111111111_1101110111010010_0010000111000000"; -- -0.13351239264011383
	pesos_i(5116) := b"0000000000000000_0000000000000000_0011010001010101_1100001111000000"; -- 0.20443366467952728
	pesos_i(5117) := b"1111111111111111_1111111111111111_1110000000110100_1100100100100000"; -- -0.12419455498456955
	pesos_i(5118) := b"1111111111111111_1111111111111111_1111000111000011_0101101010000000"; -- -0.05561289191246033
	pesos_i(5119) := b"1111111111111111_1111111111111111_1101000010010011_1100101100000000"; -- -0.1852448582649231
	pesos_i(5120) := b"0000000000000000_0000000000000000_0001110011010100_0010100110100000"; -- 0.11261234432458878
	pesos_i(5121) := b"0000000000000000_0000000000000000_0100011111111111_0000100000000000"; -- 0.2812352180480957
	pesos_i(5122) := b"0000000000000000_0000000000000000_0000110000000011_1011000000010000"; -- 0.04693127050995827
	pesos_i(5123) := b"1111111111111111_1111111111111111_1100111111100001_1100101111000000"; -- -0.18796087801456451
	pesos_i(5124) := b"0000000000000000_0000000000000000_0100001010011111_0110110010000000"; -- 0.26024511456489563
	pesos_i(5125) := b"1111111111111111_1111111111111111_1101111111001111_0110100101000000"; -- -0.1257414072751999
	pesos_i(5126) := b"0000000000000000_0000000000000000_0011001011110001_0111110100000000"; -- 0.19899731874465942
	pesos_i(5127) := b"0000000000000000_0000000000000000_0000100001110010_0111010000100000"; -- 0.03299642354249954
	pesos_i(5128) := b"1111111111111111_1111111111111111_1111000001010110_0100111111010000"; -- -0.061182986944913864
	pesos_i(5129) := b"1111111111111111_1111111111111111_1100101010101110_0100100101000000"; -- -0.2082781046628952
	pesos_i(5130) := b"0000000000000000_0000000000000000_0001101011010000_0101111001100000"; -- 0.10474195331335068
	pesos_i(5131) := b"0000000000000000_0000000000000000_0011011001100001_1101111011000000"; -- 0.21243087947368622
	pesos_i(5132) := b"1111111111111111_1111111111111111_1111001000001100_1101000000100000"; -- -0.05449198931455612
	pesos_i(5133) := b"1111111111111111_1111111111111111_1101110000001011_1000000110000000"; -- -0.1404494345188141
	pesos_i(5134) := b"0000000000000000_0000000000000000_0000110110010111_0001000010010000"; -- 0.05308631435036659
	pesos_i(5135) := b"1111111111111111_1111111111111111_1111101010000001_0101011010101000"; -- -0.021463951095938683
	pesos_i(5136) := b"1111111111111111_1111111111111111_1111011111011000_1110110100010000"; -- -0.031846221536397934
	pesos_i(5137) := b"0000000000000000_0000000000000000_0001110111001001_1110011101100000"; -- 0.1163620576262474
	pesos_i(5138) := b"1111111111111111_1111111111111111_1111111111111001_1011010001000101"; -- -9.606652020011097e-05
	pesos_i(5139) := b"1111111111111111_1111111111111111_1100010100110100_0010011000000000"; -- -0.22967302799224854
	pesos_i(5140) := b"0000000000000000_0000000000000000_0000000100110001_1011100001100000"; -- 0.004664920270442963
	pesos_i(5141) := b"0000000000000000_0000000000000000_0001111100100101_1011100011000000"; -- 0.12166933715343475
	pesos_i(5142) := b"0000000000000000_0000000000000000_0010000111110000_1100110110000000"; -- 0.13258060812950134
	pesos_i(5143) := b"1111111111111111_1111111111111111_1100101010100001_0000001011000000"; -- -0.20848067104816437
	pesos_i(5144) := b"0000000000000000_0000000000000000_0010001011000111_1000110100000000"; -- 0.13585740327835083
	pesos_i(5145) := b"1111111111111111_1111111111111111_1010011111100010_0111101100000000"; -- -0.3442004323005676
	pesos_i(5146) := b"0000000000000000_0000000000000000_0100111110010101_0111111110000000"; -- 0.31087490916252136
	pesos_i(5147) := b"1111111111111111_1111111111111111_1111000110110100_0010000001010000"; -- -0.055845241993665695
	pesos_i(5148) := b"0000000000000000_0000000000000000_0100000011010110_0100100100000000"; -- 0.2532697319984436
	pesos_i(5149) := b"1111111111111111_1111111111111111_1011010001100101_0000101010000000"; -- -0.29533323645591736
	pesos_i(5150) := b"0000000000000000_0000000000000000_0101110101110001_1010100110000000"; -- 0.36501559615135193
	pesos_i(5151) := b"1111111111111111_1111111111111111_1101000010110001_0101101000000000"; -- -0.18479382991790771
	pesos_i(5152) := b"0000000000000000_0000000000000000_0001010001111010_0011000100000000"; -- 0.079989492893219
	pesos_i(5153) := b"0000000000000000_0000000000000000_0011010111010001_1010111110000000"; -- 0.21023079752922058
	pesos_i(5154) := b"0000000000000000_0000000000000000_0010011111111110_1101111001000000"; -- 0.15623272955417633
	pesos_i(5155) := b"1111111111111111_1111111111111111_1110001001000010_0011000001000000"; -- -0.11617754399776459
	pesos_i(5156) := b"0000000000000000_0000000000000000_0010101000010010_0010101011000000"; -- 0.16433970630168915
	pesos_i(5157) := b"0000000000000000_0000000000000000_0010111011100011_1011001100000000"; -- 0.1831619143486023
	pesos_i(5158) := b"1111111111111111_1111111111111111_1101010101100011_1111010000000000"; -- -0.1664435863494873
	pesos_i(5159) := b"0000000000000000_0000000000000000_0000100101000000_1000010010110000"; -- 0.036140721291303635
	pesos_i(5160) := b"0000000000000000_0000000000000000_0010101101100000_1010101010000000"; -- 0.1694437563419342
	pesos_i(5161) := b"1111111111111111_1111111111111111_1110000111000001_1001110001000000"; -- -0.11813949048519135
	pesos_i(5162) := b"1111111111111111_1111111111111111_1011100000010111_1101110110000000"; -- -0.28088584542274475
	pesos_i(5163) := b"1111111111111111_1111111111111111_1110011100011000_1101001110000000"; -- -0.09727743268013
	pesos_i(5164) := b"1111111111111111_1111111111111111_1111010110100100_1101111001010000"; -- -0.04045305773615837
	pesos_i(5165) := b"0000000000000000_0000000000000000_0001010011110111_0011110011100000"; -- 0.0818975493311882
	pesos_i(5166) := b"0000000000000000_0000000000000000_0001111101110111_1100001110000000"; -- 0.12292119860649109
	pesos_i(5167) := b"0000000000000000_0000000000000000_0001000110100010_1000110000000000"; -- 0.06888651847839355
	pesos_i(5168) := b"1111111111111111_1111111111111111_1111110001011010_0011100010101100"; -- -0.01424833107739687
	pesos_i(5169) := b"1111111111111111_1111111111111111_1111100111111000_0111110100001000"; -- -0.023552117869257927
	pesos_i(5170) := b"1111111111111111_1111111111111111_1111101011010111_0010100000001000"; -- -0.020154474303126335
	pesos_i(5171) := b"0000000000000000_0000000000000000_0010101101110001_1100000011000000"; -- 0.16970448195934296
	pesos_i(5172) := b"0000000000000000_0000000000000000_0001110110010110_0001010001000000"; -- 0.1155712753534317
	pesos_i(5173) := b"1111111111111111_1111111111111111_1111110111101110_0000101111000000"; -- -0.00808645784854889
	pesos_i(5174) := b"0000000000000000_0000000000000000_0000100010110010_0001001111010000"; -- 0.03396724537014961
	pesos_i(5175) := b"0000000000000000_0000000000000000_0010001100101111_1001010110000000"; -- 0.13744482398033142
	pesos_i(5176) := b"1111111111111111_1111111111111111_1111011111000111_0011110101010000"; -- -0.03211609646677971
	pesos_i(5177) := b"0000000000000000_0000000000000000_0010000000000000_1100001001000000"; -- 0.12501157820224762
	pesos_i(5178) := b"1111111111111111_1111111111111111_1000101101001011_0101111010000000"; -- -0.4558812081813812
	pesos_i(5179) := b"0000000000000000_0000000000000000_0100001010001111_1101000000000000"; -- 0.2600069046020508
	pesos_i(5180) := b"0000000000000000_0000000000000000_0010110000111100_0101010001000000"; -- 0.17279554903507233
	pesos_i(5181) := b"1111111111111111_1111111111111111_1100110110100110_0010100100000000"; -- -0.1966833472251892
	pesos_i(5182) := b"0000000000000000_0000000000000000_0000101001100001_1111010111000000"; -- 0.04055725038051605
	pesos_i(5183) := b"1111111111111111_1111111111111111_1110100011010110_0101100110000000"; -- -0.0904792845249176
	pesos_i(5184) := b"0000000000000000_0000000000000000_0000101101100110_0001101110000000"; -- 0.04452678561210632
	pesos_i(5185) := b"0000000000000000_0000000000000000_0001000100001111_1100001001100000"; -- 0.06664671748876572
	pesos_i(5186) := b"0000000000000000_0000000000000000_0010111000100001_0110111001000000"; -- 0.180197611451149
	pesos_i(5187) := b"0000000000000000_0000000000000000_0001000011111000_1011011001100000"; -- 0.06629505008459091
	pesos_i(5188) := b"0000000000000000_0000000000000000_0011011110011110_0101000101000000"; -- 0.217259481549263
	pesos_i(5189) := b"0000000000000000_0000000000000000_0011001100111011_0000001110000000"; -- 0.2001192271709442
	pesos_i(5190) := b"1111111111111111_1111111111111111_1010110001111101_0010001000000000"; -- -0.32621562480926514
	pesos_i(5191) := b"0000000000000000_0000000000000000_0000001001100011_0100100010111000"; -- 0.00932745449244976
	pesos_i(5192) := b"0000000000000000_0000000000000000_0001010100000001_1011001000000000"; -- 0.08205711841583252
	pesos_i(5193) := b"1111111111111111_1111111111111111_1111010100001100_0000001110010000"; -- -0.04278543218970299
	pesos_i(5194) := b"0000000000000000_0000000000000000_0000011111101111_0000000101001000"; -- 0.03099067695438862
	pesos_i(5195) := b"0000000000000000_0000000000000000_0000100001101110_0100010111110000"; -- 0.03293263539671898
	pesos_i(5196) := b"1111111111111111_1111111111111111_1001101111101001_1001101110000000"; -- -0.3909666836261749
	pesos_i(5197) := b"1111111111111111_1111111111111111_1111010000101010_1111011000010000"; -- -0.046219464391469955
	pesos_i(5198) := b"0000000000000000_0000000000000000_0001010010111001_1101100000100000"; -- 0.08096075803041458
	pesos_i(5199) := b"0000000000000000_0000000000000000_0001101000011010_1010100111000000"; -- 0.10196934640407562
	pesos_i(5200) := b"0000000000000000_0000000000000000_0010010001110110_0110000011000000"; -- 0.14243130385875702
	pesos_i(5201) := b"0000000000000000_0000000000000000_0010100010000101_1111110000000000"; -- 0.1582944393157959
	pesos_i(5202) := b"1111111111111111_1111111111111111_1100100011010100_1111000010000000"; -- -0.21550080180168152
	pesos_i(5203) := b"0000000000000000_0000000000000000_0000001110101001_1001010111100000"; -- 0.014306418597698212
	pesos_i(5204) := b"0000000000000000_0000000000000000_0010111110110011_1100011011000000"; -- 0.1863369196653366
	pesos_i(5205) := b"0000000000000000_0000000000000000_0010001010010101_1110100001000000"; -- 0.13509990274906158
	pesos_i(5206) := b"0000000000000000_0000000000000000_0011000001100001_1110010101000000"; -- 0.18899376690387726
	pesos_i(5207) := b"1111111111111111_1111111111111111_1110000000011101_0110101110000000"; -- -0.12455108761787415
	pesos_i(5208) := b"1111111111111111_1111111111111111_1111111001110010_1101101001111100"; -- -0.006059975363314152
	pesos_i(5209) := b"0000000000000000_0000000000000000_0011000100000010_1011010000000000"; -- 0.19144749641418457
	pesos_i(5210) := b"1111111111111111_1111111111111111_1111110000100110_1100100110001100"; -- -0.015033152885735035
	pesos_i(5211) := b"0000000000000000_0000000000000000_0000001010001010_0001001011110000"; -- 0.009919341653585434
	pesos_i(5212) := b"1111111111111111_1111111111111111_1011100110011011_1010001100000000"; -- -0.2749689221382141
	pesos_i(5213) := b"1111111111111111_1111111111111111_1011001001111000_0011010100000000"; -- -0.3028532862663269
	pesos_i(5214) := b"1111111111111111_1111111111111111_1110101101000100_1001110101000000"; -- -0.08098427951335907
	pesos_i(5215) := b"1111111111111111_1111111111111111_1110100111011111_1010100110000000"; -- -0.08643093705177307
	pesos_i(5216) := b"0000000000000000_0000000000000000_0000110010001110_0001011000000000"; -- 0.04904305934906006
	pesos_i(5217) := b"0000000000000000_0000000000000000_0000010001000010_1001011100011000"; -- 0.01664108596742153
	pesos_i(5218) := b"0000000000000000_0000000000000000_0010100011110011_0101011001000000"; -- 0.15996302664279938
	pesos_i(5219) := b"0000000000000000_0000000000000000_0011100011001010_0101011000000000"; -- 0.22183740139007568
	pesos_i(5220) := b"0000000000000000_0000000000000000_0000101101110000_1011001000110000"; -- 0.044688355177640915
	pesos_i(5221) := b"0000000000000000_0000000000000000_0000001000001110_0011001111111100"; -- 0.008029221557080746
	pesos_i(5222) := b"0000000000000000_0000000000000000_0011010010000000_1010111011000000"; -- 0.2050885409116745
	pesos_i(5223) := b"0000000000000000_0000000000000000_0001110110101001_0010010111000000"; -- 0.11586223542690277
	pesos_i(5224) := b"1111111111111111_1111111111111111_1010011010101111_1001010110000000"; -- -0.3488833010196686
	pesos_i(5225) := b"1111111111111111_1111111111111111_1101110110010001_1010011111000000"; -- -0.13449622690677643
	pesos_i(5226) := b"0000000000000000_0000000000000000_0001100111101100_1000001110100000"; -- 0.10126516968011856
	pesos_i(5227) := b"0000000000000000_0000000000000000_0010000000111011_1111011110000000"; -- 0.1259150207042694
	pesos_i(5228) := b"0000000000000000_0000000000000000_0010100000110011_0001100100000000"; -- 0.15702968835830688
	pesos_i(5229) := b"0000000000000000_0000000000000000_0010000010001000_1100111100000000"; -- 0.1270875334739685
	pesos_i(5230) := b"1111111111111111_1111111111111111_1100010100110100_1001100011000000"; -- -0.22966618835926056
	pesos_i(5231) := b"1111111111111111_1111111111111111_1010010000000110_1010010100000000"; -- -0.35927361249923706
	pesos_i(5232) := b"1111111111111111_1111111111111111_1100011111100111_1110101000000000"; -- -0.21911752223968506
	pesos_i(5233) := b"1111111111111111_1111111111111111_1110111110111011_0001111010100000"; -- -0.06355103105306625
	pesos_i(5234) := b"0000000000000000_0000000000000000_0001000011101101_1111111010000000"; -- 0.06613150238990784
	pesos_i(5235) := b"0000000000000000_0000000000000000_0011111001101001_1111001000000000"; -- 0.24380409717559814
	pesos_i(5236) := b"1111111111111111_1111111111111111_1110100000101100_1011100000000000"; -- -0.09306764602661133
	pesos_i(5237) := b"0000000000000000_0000000000000000_0000100010101000_0010110111100000"; -- 0.03381621092557907
	pesos_i(5238) := b"1111111111111111_1111111111111111_1100101101101011_1110010010000000"; -- -0.20538493990898132
	pesos_i(5239) := b"0000000000000000_0000000000000000_0101001110111011_1100011110000000"; -- 0.3270840346813202
	pesos_i(5240) := b"0000000000000000_0000000000000000_0000110101110110_1001101111000000"; -- 0.05259107053279877
	pesos_i(5241) := b"0000000000000000_0000000000000000_0001001000101000_1110100111100000"; -- 0.07093679159879684
	pesos_i(5242) := b"1111111111111111_1111111111111111_1101101001101110_0001010101000000"; -- -0.14675776660442352
	pesos_i(5243) := b"1111111111111111_1111111111111111_1011010100110000_0101000010000000"; -- -0.2922315299510956
	pesos_i(5244) := b"0000000000000000_0000000000000000_0001000001110010_1010101011000000"; -- 0.0642496794462204
	pesos_i(5245) := b"1111111111111111_1111111111111111_1111101011001011_1011101010110000"; -- -0.020328838378190994
	pesos_i(5246) := b"1111111111111111_1111111111111111_1111010100101011_1000010011010000"; -- -0.04230470582842827
	pesos_i(5247) := b"0000000000000000_0000000000000000_0001010100010001_1101010110000000"; -- 0.08230337500572205
	pesos_i(5248) := b"0000000000000000_0000000000000000_0100001011111100_1000011010000000"; -- 0.2616657316684723
	pesos_i(5249) := b"1111111111111111_1111111111111111_1011100100100011_0011101100000000"; -- -0.27680617570877075
	pesos_i(5250) := b"0000000000000000_0000000000000000_0001101001011011_0110101100000000"; -- 0.10295742750167847
	pesos_i(5251) := b"1111111111111111_1111111111111111_1101110011010000_0010011110000000"; -- -0.13744881749153137
	pesos_i(5252) := b"0000000000000000_0000000000000000_0010010010001100_1010111001000000"; -- 0.1427716165781021
	pesos_i(5253) := b"0000000000000000_0000000000000000_0000010000111111_1010000110010000"; -- 0.016595933586359024
	pesos_i(5254) := b"0000000000000000_0000000000000000_0100101001010010_0100101100000000"; -- 0.29031819105148315
	pesos_i(5255) := b"0000000000000000_0000000000000000_0001000111101100_1011111111100000"; -- 0.07001876085996628
	pesos_i(5256) := b"1111111111111111_1111111111111111_1010000001110101_0000111100000000"; -- -0.37321382761001587
	pesos_i(5257) := b"0000000000000000_0000000000000000_0001110001101110_1100110010000000"; -- 0.11106565594673157
	pesos_i(5258) := b"0000000000000000_0000000000000000_0001111001111011_1110010100100000"; -- 0.11907798796892166
	pesos_i(5259) := b"0000000000000000_0000000000000000_0000110001100101_1111110101010000"; -- 0.048431236296892166
	pesos_i(5260) := b"1111111111111111_1111111111111111_1100111101001000_1010001110000000"; -- -0.19029787182807922
	pesos_i(5261) := b"1111111111111111_1111111111111111_1111001011101010_1100100101110000"; -- -0.05110493674874306
	pesos_i(5262) := b"0000000000000000_0000000000000000_0000110010111110_0110000100110000"; -- 0.04977996274828911
	pesos_i(5263) := b"0000000000000000_0000000000000000_0000010000101101_0010110101010000"; -- 0.016314346343278885
	pesos_i(5264) := b"0000000000000000_0000000000000000_0000011011100010_0010011111001000"; -- 0.02688835747539997
	pesos_i(5265) := b"1111111111111111_1111111111111111_1111011010010100_0111011010010000"; -- -0.03679713234305382
	pesos_i(5266) := b"0000000000000000_0000000000000000_0001101001010101_1011001010000000"; -- 0.10287013649940491
	pesos_i(5267) := b"1111111111111111_1111111111111111_1110000111000010_0011010100100000"; -- -0.11813037842512131
	pesos_i(5268) := b"1111111111111111_1111111111111111_1111100101100100_0101010110001000"; -- -0.025812773033976555
	pesos_i(5269) := b"1111111111111111_1111111111111111_1111011010010000_1100010111110000"; -- -0.03685343638062477
	pesos_i(5270) := b"1111111111111111_1111111111111111_1001101110001100_0111011100000000"; -- -0.39238792657852173
	pesos_i(5271) := b"0000000000000000_0000000000000000_0000101010110000_1010000100010000"; -- 0.041757646948099136
	pesos_i(5272) := b"0000000000000000_0000000000000000_0001100001010101_0000101110100000"; -- 0.09504768997430801
	pesos_i(5273) := b"1111111111111111_1111111111111111_1100110101100111_0111011011000000"; -- -0.19764001667499542
	pesos_i(5274) := b"0000000000000000_0000000000000000_0010000000111001_1011111111000000"; -- 0.12588118016719818
	pesos_i(5275) := b"1111111111111111_1111111111111111_1110010101101001_1000010100100000"; -- -0.10385864228010178
	pesos_i(5276) := b"0000000000000000_0000000000000000_0001001111110011_1111011011000000"; -- 0.07794134318828583
	pesos_i(5277) := b"1111111111111111_1111111111111111_1111010001011101_1001110110010000"; -- -0.04544654116034508
	pesos_i(5278) := b"1111111111111111_1111111111111111_1111111010010101_0100011010001100"; -- -0.005534735508263111
	pesos_i(5279) := b"1111111111111111_1111111111111111_1101011000001100_0110111011000000"; -- -0.16387279331684113
	pesos_i(5280) := b"1111111111111111_1111111111111111_1101001001101000_0001110011000000"; -- -0.1780988723039627
	pesos_i(5281) := b"0000000000000000_0000000000000000_0011010011001000_1010101000000000"; -- 0.20618689060211182
	pesos_i(5282) := b"0000000000000000_0000000000000000_0011010001100000_0101010001000000"; -- 0.20459486544132233
	pesos_i(5283) := b"1111111111111111_1111111111111111_1110000100000011_0111000010100000"; -- -0.12104126065969467
	pesos_i(5284) := b"0000000000000000_0000000000000000_0100000101010111_0101000100000000"; -- 0.2552385926246643
	pesos_i(5285) := b"0000000000000000_0000000000000000_0000001111001111_1110011001001100"; -- 0.014891046099364758
	pesos_i(5286) := b"0000000000000000_0000000000000000_0010110010000110_0111111111000000"; -- 0.17392729222774506
	pesos_i(5287) := b"1111111111111111_1111111111111111_1110011111000010_0111110001100000"; -- -0.09468863159418106
	pesos_i(5288) := b"0000000000000000_0000000000000000_0000001100001010_1010101010110100"; -- 0.011881512589752674
	pesos_i(5289) := b"1111111111111111_1111111111111111_1101101100011110_1100111101000000"; -- -0.1440611332654953
	pesos_i(5290) := b"1111111111111111_1111111111111111_1110111111001111_0000101101100000"; -- -0.06324700266122818
	pesos_i(5291) := b"0000000000000000_0000000000000000_0001011010110101_1100001111100000"; -- 0.08871101588010788
	pesos_i(5292) := b"1111111111111111_1111111111111111_1100000001000011_0001101100000000"; -- -0.24897605180740356
	pesos_i(5293) := b"1111111111111111_1111111111111111_1111010101110100_0110111001100000"; -- -0.041192151606082916
	pesos_i(5294) := b"1111111111111111_1111111111111111_1001001111100101_1011100110000000"; -- -0.42227593064308167
	pesos_i(5295) := b"1111111111111111_1111111111111111_1101010101110100_0100000000000000"; -- -0.16619491577148438
	pesos_i(5296) := b"0000000000000000_0000000000000000_0011011100110110_0100000111000000"; -- 0.21567164361476898
	pesos_i(5297) := b"1111111111111111_1111111111111111_1010101001110011_1001000100000000"; -- -0.33417409658432007
	pesos_i(5298) := b"1111111111111111_1111111111111111_1101010110111111_0111111100000000"; -- -0.16504675149917603
	pesos_i(5299) := b"0000000000000000_0000000000000000_0001010011000011_0100111011000000"; -- 0.08110515773296356
	pesos_i(5300) := b"0000000000000000_0000000000000000_0010110010000011_0110001001000000"; -- 0.17387975752353668
	pesos_i(5301) := b"1111111111111111_1111111111111111_1110001001011011_1011101000000000"; -- -0.11578786373138428
	pesos_i(5302) := b"1111111111111111_1111111111111111_1111101111011101_1001010010001000"; -- -0.016150204464793205
	pesos_i(5303) := b"0000000000000000_0000000000000000_0000111100101111_0111111000010000"; -- 0.0593184269964695
	pesos_i(5304) := b"1111111111111111_1111111111111111_1010110110001110_0000011000000000"; -- -0.32205164432525635
	pesos_i(5305) := b"1111111111111111_1111111111111111_1111001111011110_0011111111000000"; -- -0.04738999903202057
	pesos_i(5306) := b"1111111111111111_1111111111111111_1100101101010010_1001110000000000"; -- -0.20577073097229004
	pesos_i(5307) := b"0000000000000000_0000000000000000_0010000011001000_0000111110000000"; -- 0.12805268168449402
	pesos_i(5308) := b"0000000000000000_0000000000000000_0000000100111110_0101011101001100"; -- 0.004857498221099377
	pesos_i(5309) := b"1111111111111111_1111111111111111_1111001111001101_0110000001010000"; -- -0.04764745756983757
	pesos_i(5310) := b"0000000000000000_0000000000000000_0010101000011100_0011011110000000"; -- 0.16449305415153503
	pesos_i(5311) := b"1111111111111111_1111111111111111_1101000010111100_1000111110000000"; -- -0.18462279438972473
	pesos_i(5312) := b"0000000000000000_0000000000000000_0010000011001100_0100111111000000"; -- 0.12811754643917084
	pesos_i(5313) := b"0000000000000000_0000000000000000_0010100101011001_0111010000000000"; -- 0.16152119636535645
	pesos_i(5314) := b"1111111111111111_1111111111111111_1111000011100110_1001000111110000"; -- -0.05898177996277809
	pesos_i(5315) := b"0000000000000000_0000000000000000_0000100011010110_0001111000100000"; -- 0.03451717644929886
	pesos_i(5316) := b"0000000000000000_0000000000000000_0010000010100001_0100111100000000"; -- 0.12746137380599976
	pesos_i(5317) := b"0000000000000000_0000000000000000_0010101110001111_0001110110000000"; -- 0.17015251517295837
	pesos_i(5318) := b"1111111111111111_1111111111111111_1100011010011011_1000001111000000"; -- -0.22418953478336334
	pesos_i(5319) := b"0000000000000000_0000000000000000_0010111111111111_0001000110000000"; -- 0.18748578429222107
	pesos_i(5320) := b"0000000000000000_0000000000000000_0011101111100100_1100011001000000"; -- 0.23395957052707672
	pesos_i(5321) := b"1111111111111111_1111111111111111_1111010001000010_1001110100110000"; -- -0.04585855081677437
	pesos_i(5322) := b"1111111111111111_1111111111111111_1011110100111001_1100111010000000"; -- -0.2608366906642914
	pesos_i(5323) := b"0000000000000000_0000000000000000_0010111111110110_1001111110000000"; -- 0.18735691905021667
	pesos_i(5324) := b"1111111111111111_1111111111111111_1110100001111010_0011000010000000"; -- -0.0918855369091034
	pesos_i(5325) := b"0000000000000000_0000000000000000_0010000111011010_0010011111000000"; -- 0.13223503530025482
	pesos_i(5326) := b"0000000000000000_0000000000000000_0101110101001010_0010110010000000"; -- 0.3644130527973175
	pesos_i(5327) := b"0000000000000000_0000000000000000_0001010001010000_1010110111100000"; -- 0.07935606688261032
	pesos_i(5328) := b"0000000000000000_0000000000000000_0001000000010100_1010101001100000"; -- 0.06281533092260361
	pesos_i(5329) := b"0000000000000000_0000000000000000_0011001101010101_0010010110000000"; -- 0.20051798224449158
	pesos_i(5330) := b"1111111111111111_1111111111111111_1101011111000111_0101110101000000"; -- -0.1571141928434372
	pesos_i(5331) := b"0000000000000000_0000000000000000_0001101100000000_1011111001100000"; -- 0.10548009723424911
	pesos_i(5332) := b"1111111111111111_1111111111111111_1101000011101010_0011111110000000"; -- -0.18392565846443176
	pesos_i(5333) := b"0000000000000000_0000000000000000_0011111110101111_0110011110000000"; -- 0.24877020716667175
	pesos_i(5334) := b"0000000000000000_0000000000000000_0000110100111100_0001100100110000"; -- 0.05169827863574028
	pesos_i(5335) := b"1111111111111111_1111111111111111_1011010111011111_1001010100000000"; -- -0.28955715894699097
	pesos_i(5336) := b"1111111111111111_1111111111111111_1011010110000100_0011001100000000"; -- -0.29095155000686646
	pesos_i(5337) := b"0000000000000000_0000000000000000_0011110010011000_1000101001000000"; -- 0.2367025762796402
	pesos_i(5338) := b"1111111111111111_1111111111111111_1110011011010110_1010011111100000"; -- -0.09828711301088333
	pesos_i(5339) := b"1111111111111111_1111111111111111_1110011101011001_1101100010000000"; -- -0.09628531336784363
	pesos_i(5340) := b"1111111111111111_1111111111111111_1011111100011101_1111010110000000"; -- -0.25344911217689514
	pesos_i(5341) := b"0000000000000000_0000000000000000_0000101100011110_0101100100000000"; -- 0.04343181848526001
	pesos_i(5342) := b"1111111111111111_1111111111111111_1101111111100111_0010000110000000"; -- -0.12537947297096252
	pesos_i(5343) := b"1111111111111111_1111111111111111_1110111100010100_0011010101000000"; -- -0.06609790027141571
	pesos_i(5344) := b"0000000000000000_0000000000000000_0010100100001101_1101110110000000"; -- 0.16036781668663025
	pesos_i(5345) := b"0000000000000000_0000000000000000_0001110110010011_0111000000100000"; -- 0.11553097516298294
	pesos_i(5346) := b"0000000000000000_0000000000000000_0011001111111010_0110000110000000"; -- 0.2030392587184906
	pesos_i(5347) := b"0000000000000000_0000000000000000_0010100011001100_0111101111000000"; -- 0.15937016904354095
	pesos_i(5348) := b"0000000000000000_0000000000000000_0010001001111101_0001000010000000"; -- 0.1347208321094513
	pesos_i(5349) := b"0000000000000000_0000000000000000_0010100101110000_0100100011000000"; -- 0.1618695706129074
	pesos_i(5350) := b"0000000000000000_0000000000000000_0011101101010000_1001011101000000"; -- 0.23169846832752228
	pesos_i(5351) := b"0000000000000000_0000000000000000_0100000000011010_0101110000000000"; -- 0.25040221214294434
	pesos_i(5352) := b"0000000000000000_0000000000000000_0010000000000010_1100011000000000"; -- 0.12504231929779053
	pesos_i(5353) := b"1111111111111111_1111111111111111_1100000110110111_0110001111000000"; -- -0.24329544603824615
	pesos_i(5354) := b"1111111111111111_1111111111111111_0101011100100111_0101010100000000"; -- -0.6595560908317566
	pesos_i(5355) := b"0000000000000000_0000000000000000_0100000011010011_0111110100000000"; -- 0.2532270550727844
	pesos_i(5356) := b"0000000000000000_0000000000000000_0011101111101011_1111001101000000"; -- 0.2340690642595291
	pesos_i(5357) := b"0000000000000000_0000000000000000_0010111011011101_1010010001000000"; -- 0.18306948244571686
	pesos_i(5358) := b"0000000000000000_0000000000000000_0001001000110100_1001111110000000"; -- 0.07111546397209167
	pesos_i(5359) := b"1111111111111111_1111111111111111_0110011001101110_0100001100000000"; -- -0.599880039691925
	pesos_i(5360) := b"1111111111111111_1111111111111111_1100000011101101_0000011100000000"; -- -0.24638324975967407
	pesos_i(5361) := b"0000000000000000_0000000000000000_0001101000110111_1001010100000000"; -- 0.10241061449050903
	pesos_i(5362) := b"0000000000000000_0000000000000000_0000101100010000_0111110000110000"; -- 0.043220292776823044
	pesos_i(5363) := b"0000000000000000_0000000000000000_0000110110111101_1011110110010000"; -- 0.053676459938287735
	pesos_i(5364) := b"1111111111111111_1111111111111111_1101010010000011_0000000011000000"; -- -0.16987605392932892
	pesos_i(5365) := b"0000000000000000_0000000000000000_0010000010000111_1100110001000000"; -- 0.12707211077213287
	pesos_i(5366) := b"1111111111111111_1111111111111111_1111110110000001_1110101001111100"; -- -0.009736389853060246
	pesos_i(5367) := b"0000000000000000_0000000000000000_0100011110110101_1000001010000000"; -- 0.2801133692264557
	pesos_i(5368) := b"1111111111111111_1111111111111111_1111101100001111_1010100011101000"; -- -0.019292300567030907
	pesos_i(5369) := b"1111111111111111_1111111111111111_1111001010010101_1111010101000000"; -- -0.052399322390556335
	pesos_i(5370) := b"1111111111111111_1111111111111111_1011100010100001_1100110010000000"; -- -0.27878114581108093
	pesos_i(5371) := b"1111111111111111_1111111111111111_1011011011001000_0000000110000000"; -- -0.28601065278053284
	pesos_i(5372) := b"1111111111111111_1111111111111111_1110111001100011_0101101011000000"; -- -0.06879647076129913
	pesos_i(5373) := b"0000000000000000_0000000000000000_0001101011001111_1000010000000000"; -- 0.10472893714904785
	pesos_i(5374) := b"1111111111111111_1111111111111111_1101010010000110_0000101110000000"; -- -0.16982963681221008
	pesos_i(5375) := b"0000000000000000_0000000000000000_0001100011010111_1101110011100000"; -- 0.09704380482435226
	pesos_i(5376) := b"0000000000000000_0000000000000000_0100011011100001_1110000100000000"; -- 0.27688413858413696
	pesos_i(5377) := b"1111111111111111_1111111111111111_1001000110110111_1011100010000000"; -- -0.43079039454460144
	pesos_i(5378) := b"0000000000000000_0000000000000000_0001100001101010_0110000100100000"; -- 0.09537322074174881
	pesos_i(5379) := b"0000000000000000_0000000000000000_0010011101011001_1110001001000000"; -- 0.15371526777744293
	pesos_i(5380) := b"1111111111111111_1111111111111111_1100000011010001_1111010111000000"; -- -0.24679626524448395
	pesos_i(5381) := b"0000000000000000_0000000000000000_0100000001100111_1010010100000000"; -- 0.25158149003982544
	pesos_i(5382) := b"0000000000000000_0000000000000000_0111100001100000_1000110010000000"; -- 0.47022321820259094
	pesos_i(5383) := b"0000000000000000_0000000000000000_0001000000111110_1101111101100000"; -- 0.0634593591094017
	pesos_i(5384) := b"1111111111111111_1111111111111111_1000111110011010_0011010010000000"; -- -0.4390532672405243
	pesos_i(5385) := b"0000000000000000_0000000000000000_0100000011111011_1010101110000000"; -- 0.2538401782512665
	pesos_i(5386) := b"0000000000000000_0000000000000000_0010011010101001_0100011010000000"; -- 0.15102043747901917
	pesos_i(5387) := b"1111111111111111_1111111111111111_1101001000101101_1101100001000000"; -- -0.17898796498775482
	pesos_i(5388) := b"1111111111111111_1111111111111111_1110010111100111_1110110011100000"; -- -0.10192985087633133
	pesos_i(5389) := b"0000000000000000_0000000000000000_0001010101001110_0111111100100000"; -- 0.08322901278734207
	pesos_i(5390) := b"0000000000000000_0000000000000000_0011001101000111_0001100100000000"; -- 0.20030361413955688
	pesos_i(5391) := b"1111111111111111_1111111111111111_1101000101111100_1101011000000000"; -- -0.18168890476226807
	pesos_i(5392) := b"1111111111111111_1111111111111111_1111000011110101_1001000000100000"; -- -0.05875300616025925
	pesos_i(5393) := b"0000000000000000_0000000000000000_0101011011011010_1100101000000000"; -- 0.33927595615386963
	pesos_i(5394) := b"0000000000000000_0000000000000000_0101011011110110_0110001010000000"; -- 0.3396970331668854
	pesos_i(5395) := b"0000000000000000_0000000000000000_0011110100001011_0000100000000000"; -- 0.2384495735168457
	pesos_i(5396) := b"0000000000000000_0000000000000000_0101000100100010_1000000100000000"; -- 0.316932737827301
	pesos_i(5397) := b"1111111111111111_1111111111111111_1101011101111010_1000010111000000"; -- -0.1582867056131363
	pesos_i(5398) := b"1111111111111111_1111111111111111_0110010111010011_1001111000000000"; -- -0.602239727973938
	pesos_i(5399) := b"1111111111111111_1111111111111111_1100110100000010_0100011001000000"; -- -0.19918404519557953
	pesos_i(5400) := b"1111111111111111_1111111111111111_1011010110110101_0010111110000000"; -- -0.29020407795906067
	pesos_i(5401) := b"1111111111111111_1111111111111111_1110101011100101_1010010101100000"; -- -0.08243338018655777
	pesos_i(5402) := b"1111111111111111_1111111111111111_1110000111101101_0011010011100000"; -- -0.117474265396595
	pesos_i(5403) := b"0000000000000000_0000000000000000_0010100111100001_1001101111000000"; -- 0.16359876096248627
	pesos_i(5404) := b"1111111111111111_1111111111111111_1100110100011000_0100101000000000"; -- -0.19884812831878662
	pesos_i(5405) := b"0000000000000000_0000000000000000_0101100011001001_1100011000000000"; -- 0.346828818321228
	pesos_i(5406) := b"1111111111111111_1111111111111111_1111000000101100_1001100100000000"; -- -0.061819493770599365
	pesos_i(5407) := b"0000000000000000_0000000000000000_0100000111010111_0101101110000000"; -- 0.25719234347343445
	pesos_i(5408) := b"1111111111111111_1111111111111111_1101001011011111_1110011100000000"; -- -0.17627102136611938
	pesos_i(5409) := b"0000000000000000_0000000000000000_0100110101110100_1100111010000000"; -- 0.3025635778903961
	pesos_i(5410) := b"0000000000000000_0000000000000000_0101010000101000_0100101100000000"; -- 0.32873982191085815
	pesos_i(5411) := b"0000000000000000_0000000000000000_0011000111001100_0110001100000000"; -- 0.19452494382858276
	pesos_i(5412) := b"0000000000000000_0000000000000000_0001000000101110_1000100100100000"; -- 0.06321007758378983
	pesos_i(5413) := b"0000000000000000_0000000000000000_0001000111001001_1010000111000000"; -- 0.06948290765285492
	pesos_i(5414) := b"0000000000000000_0000000000000000_0010011001000100_1100010001000000"; -- 0.14948679506778717
	pesos_i(5415) := b"0000000000000000_0000000000000000_0011001001011011_0001010001000000"; -- 0.1967022567987442
	pesos_i(5416) := b"1111111111111111_1111111111111111_1101000000011100_1111011010000000"; -- -0.18705806136131287
	pesos_i(5417) := b"0000000000000000_0000000000000000_0011111000100010_0001000100000000"; -- 0.24270731210708618
	pesos_i(5418) := b"0000000000000000_0000000000000000_0010000000110100_0110100101000000"; -- 0.1257997304201126
	pesos_i(5419) := b"1111111111111111_1111111111111111_1001010101111011_1010001010000000"; -- -0.4160822331905365
	pesos_i(5420) := b"1111111111111111_1111111111111111_1110001101100100_1010000100100000"; -- -0.11174576729536057
	pesos_i(5421) := b"0000000000000000_0000000000000000_0110101001001111_0001111110000000"; -- 0.4152698218822479
	pesos_i(5422) := b"1111111111111111_1111111111111111_0110110011101011_1101111100000000"; -- -0.5745258927345276
	pesos_i(5423) := b"0000000000000000_0000000000000000_0010110011101011_1011010001000000"; -- 0.17547155916690826
	pesos_i(5424) := b"1111111111111111_1111111111111111_1111000001001111_0110010111110000"; -- -0.06128847971558571
	pesos_i(5425) := b"1111111111111111_1111111111111111_1110110110110011_1001010001100000"; -- -0.07147858291864395
	pesos_i(5426) := b"1111111111111111_1111111111111111_0111101100110110_1001101000000000"; -- -0.5186980962753296
	pesos_i(5427) := b"1111111111111111_1111111111111111_1110011101010011_1111111101000000"; -- -0.09637455642223358
	pesos_i(5428) := b"0000000000000000_0000000000000000_0010101101011100_1100001011000000"; -- 0.16938416659832
	pesos_i(5429) := b"1111111111111111_1111111111111111_1010100000010011_1001011010000000"; -- -0.3434511125087738
	pesos_i(5430) := b"0000000000000000_0000000000000000_0100001001100000_0100011010000000"; -- 0.25928154587745667
	pesos_i(5431) := b"1111111111111111_1111111111111111_1100110110011101_1110000011000000"; -- -0.19680972397327423
	pesos_i(5432) := b"1111111111111111_1111111111111111_1001110111111100_0100101010000000"; -- -0.38286909461021423
	pesos_i(5433) := b"1111111111111111_1111111111111111_1101001011001000_0001000110000000"; -- -0.17663469910621643
	pesos_i(5434) := b"0000000000000000_0000000000000000_0000011011010100_1100100000001000"; -- 0.026684286072850227
	pesos_i(5435) := b"0000000000000000_0000000000000000_0011011000011111_0100010101000000"; -- 0.2114146500825882
	pesos_i(5436) := b"1111111111111111_1111111111111111_1101001110101100_0010111000000000"; -- -0.17315399646759033
	pesos_i(5437) := b"0000000000000000_0000000000000000_0100110110000110_1011010000000000"; -- 0.30283665657043457
	pesos_i(5438) := b"1111111111111111_1111111111111111_1111010100101010_0110111110000000"; -- -0.042321234941482544
	pesos_i(5439) := b"0000000000000000_0000000000000000_0010011011000000_1011010011000000"; -- 0.15137796103954315
	pesos_i(5440) := b"0000000000000000_0000000000000000_0001111011111110_0001101110100000"; -- 0.12106487900018692
	pesos_i(5441) := b"1111111111111111_1111111111111111_1100000011000001_1001010110000000"; -- -0.24704614281654358
	pesos_i(5442) := b"0000000000000000_0000000000000000_0010100111110100_0011001011000000"; -- 0.16388241946697235
	pesos_i(5443) := b"0000000000000000_0000000000000000_0011100100101000_0111010001000000"; -- 0.22327353060245514
	pesos_i(5444) := b"1111111111111111_1111111111111111_1101100111100011_0000101011000000"; -- -0.14887936413288116
	pesos_i(5445) := b"1111111111111111_1111111111111111_1111011001011111_0001100000000000"; -- -0.03761148452758789
	pesos_i(5446) := b"0000000000000000_0000000000000000_0010111110001000_0010100000000000"; -- 0.18567132949829102
	pesos_i(5447) := b"1111111111111111_1111111111111111_1110010000101000_1100111011100000"; -- -0.10875231772661209
	pesos_i(5448) := b"0000000000000000_0000000000000000_0010000011101000_1010011110000000"; -- 0.12855002284049988
	pesos_i(5449) := b"1111111111111111_1111111111111111_1111101001000101_1001011110010000"; -- -0.02237560972571373
	pesos_i(5450) := b"1111111111111111_1111111111111111_1011101010000101_1011101110000000"; -- -0.2713969051837921
	pesos_i(5451) := b"1111111111111111_1111111111111111_1101100101001000_0110101010000000"; -- -0.15123876929283142
	pesos_i(5452) := b"0000000000000000_0000000000000000_0100001001110010_1011111100000000"; -- 0.2595633864402771
	pesos_i(5453) := b"0000000000000000_0000000000000000_0001101001101001_1111111101000000"; -- 0.10317988693714142
	pesos_i(5454) := b"0000000000000000_0000000000000000_0000011100110100_0101101001001000"; -- 0.028142588213086128
	pesos_i(5455) := b"1111111111111111_1111111111111111_1010111111001100_1100110110000000"; -- -0.31328120827674866
	pesos_i(5456) := b"1111111111111111_1111111111111111_1101000010111100_0100101110000000"; -- -0.18462684750556946
	pesos_i(5457) := b"0000000000000000_0000000000000000_0001000001100001_1101100001100000"; -- 0.06399299949407578
	pesos_i(5458) := b"1111111111111111_1111111111111111_1110110101010010_1001010010100000"; -- -0.07295867055654526
	pesos_i(5459) := b"0000000000000000_0000000000000000_0011001101010001_1100011100000000"; -- 0.2004665732383728
	pesos_i(5460) := b"1111111111111111_1111111111111111_1010111100011001_1111111110000000"; -- -0.3160095512866974
	pesos_i(5461) := b"0000000000000000_0000000000000000_0001101000110010_1000001111100000"; -- 0.10233329981565475
	pesos_i(5462) := b"1111111111111111_1111111111111111_1101000010011111_0101000110000000"; -- -0.1850689947605133
	pesos_i(5463) := b"1111111111111111_1111111111111111_1001011101000100_0111110110000000"; -- -0.4091111719608307
	pesos_i(5464) := b"1111111111111111_1111111111111111_1111110111101000_1101011010001000"; -- -0.00816592387855053
	pesos_i(5465) := b"0000000000000000_0000000000000000_0001101110111111_1110001001100000"; -- 0.10839667171239853
	pesos_i(5466) := b"0000000000000000_0000000000000000_0001010101000000_0101000001000000"; -- 0.08301259577274323
	pesos_i(5467) := b"0000000000000000_0000000000000000_0000101100110010_0010101110100000"; -- 0.043734289705753326
	pesos_i(5468) := b"1111111111111111_1111111111111111_1101110000110010_1001111010000000"; -- -0.1398526132106781
	pesos_i(5469) := b"1111111111111111_1111111111111111_1111100011011101_0001111011110000"; -- -0.02787596359848976
	pesos_i(5470) := b"0000000000000000_0000000000000000_0011100001111010_0111010010000000"; -- 0.22061851620674133
	pesos_i(5471) := b"0000000000000000_0000000000000000_0001100110111011_1100011000000000"; -- 0.10052144527435303
	pesos_i(5472) := b"1111111111111111_1111111111111111_1111100110101011_1111011100100000"; -- -0.02471976727247238
	pesos_i(5473) := b"1111111111111111_1111111111111111_1100110010000010_1111000001000000"; -- -0.2011270374059677
	pesos_i(5474) := b"0000000000000000_0000000000000000_0011111110110111_0111010100000000"; -- 0.24889308214187622
	pesos_i(5475) := b"1111111111111111_1111111111111111_1101010101111111_0101100101000000"; -- -0.1660255640745163
	pesos_i(5476) := b"0000000000000000_0000000000000000_0001101000010110_0010110111100000"; -- 0.10190092772245407
	pesos_i(5477) := b"0000000000000000_0000000000000000_0010111001101010_1100011010000000"; -- 0.18131676316261292
	pesos_i(5478) := b"0000000000000000_0000000000000000_0010010011101111_1101000100000000"; -- 0.14428430795669556
	pesos_i(5479) := b"0000000000000000_0000000000000000_0000101110000111_1001101100000000"; -- 0.045037925243377686
	pesos_i(5480) := b"1111111111111111_1111111111111111_1111111000101111_0011111111010110"; -- -0.0070915319956839085
	pesos_i(5481) := b"0000000000000000_0000000000000000_0000101111101011_0001100011110000"; -- 0.046556051820516586
	pesos_i(5482) := b"1111111111111111_1111111111111110_1111000110111001_0010101000000000"; -- -1.055768370628357
	pesos_i(5483) := b"0000000000000000_0000000000000000_0111010111100101_1100100110000000"; -- 0.46053752303123474
	pesos_i(5484) := b"0000000000000000_0000000000000000_0001010111001001_0010101111100000"; -- 0.08510088175535202
	pesos_i(5485) := b"1111111111111111_1111111111111111_1111010010001110_0101110111100000"; -- -0.04470265656709671
	pesos_i(5486) := b"0000000000000000_0000000000000000_0010011000100010_1100001100000000"; -- 0.1489679217338562
	pesos_i(5487) := b"0000000000000000_0000000000000000_0001011011110011_1110110100100000"; -- 0.08965951949357986
	pesos_i(5488) := b"1111111111111111_1111111111111111_1101100110111000_1110000110000000"; -- -0.14952269196510315
	pesos_i(5489) := b"0000000000000000_0000000000000000_0001100110010000_1000001110000000"; -- 0.09986135363578796
	pesos_i(5490) := b"1111111111111111_1111111111111111_1110110011001001_0011110000100000"; -- -0.07505439966917038
	pesos_i(5491) := b"1111111111111111_1111111111111111_1011110000110011_1011100000000000"; -- -0.26483583450317383
	pesos_i(5492) := b"1111111111111111_1111111111111111_1111011011011000_0100011001100000"; -- -0.03576240688562393
	pesos_i(5493) := b"0000000000000000_0000000000000000_0001010001101010_0011000011100000"; -- 0.0797453448176384
	pesos_i(5494) := b"0000000000000000_0000000000000000_0011111101001100_1001011010000000"; -- 0.2472623884677887
	pesos_i(5495) := b"1111111111111111_1111111111111111_1110011100100111_1100110011100000"; -- -0.09704894572496414
	pesos_i(5496) := b"0000000000000000_0000000000000000_0000100000111111_0000111111000000"; -- 0.03221224248409271
	pesos_i(5497) := b"1111111111111111_1111111111111111_1101111101100001_0001011110000000"; -- -0.12742474675178528
	pesos_i(5498) := b"1111111111111111_1111111111111111_1110001111111101_0000100110000000"; -- -0.10942021012306213
	pesos_i(5499) := b"1111111111111111_1111111111111111_1100000111110011_1000011110000000"; -- -0.24237778782844543
	pesos_i(5500) := b"0000000000000000_0000000000000000_0000100101101100_0001110101010000"; -- 0.03680594637989998
	pesos_i(5501) := b"1111111111111111_1111111111111111_1010101000000111_1111101010000000"; -- -0.33581575751304626
	pesos_i(5502) := b"1111111111111111_1111111111111111_0110101001101101_1111110000000000"; -- -0.5842592716217041
	pesos_i(5503) := b"0000000000000000_0000000000000000_0011110000010010_0111111011000000"; -- 0.23465721309185028
	pesos_i(5504) := b"0000000000000000_0000000000000000_0100100101111001_1111100110000000"; -- 0.28701743483543396
	pesos_i(5505) := b"1111111111111111_1111111111111111_1001001100000110_1101110100000000"; -- -0.42567652463912964
	pesos_i(5506) := b"1111111111111111_1111111111111111_1101110011000001_1011010010000000"; -- -0.13766929507255554
	pesos_i(5507) := b"0000000000000000_0000000000000000_0100100100111101_1010000010000000"; -- 0.28609660267829895
	pesos_i(5508) := b"1111111111111111_1111111111111111_1110011001110011_0100011100000000"; -- -0.09980350732803345
	pesos_i(5509) := b"0000000000000000_0000000000000000_0011111010001010_1101110010000000"; -- 0.24430635571479797
	pesos_i(5510) := b"1111111111111111_1111111111111111_1110010110000001_1101100100000000"; -- -0.10348743200302124
	pesos_i(5511) := b"0000000000000000_0000000000000000_0101111101111011_0110110010000000"; -- 0.37297704815864563
	pesos_i(5512) := b"0000000000000000_0000000000000000_0001000111010011_1101110011000000"; -- 0.06963901221752167
	pesos_i(5513) := b"0000000000000000_0000000000000000_0000000101111100_1001001101100010"; -- 0.0058071245439350605
	pesos_i(5514) := b"1111111111111111_1111111111111111_0111101101101111_1011100000000000"; -- -0.5178265571594238
	pesos_i(5515) := b"1111111111111111_1111111111111111_1111000010101001_1000001001000000"; -- -0.059913501143455505
	pesos_i(5516) := b"0000000000000000_0000000000000000_0001101110111110_0101010000000000"; -- 0.10837292671203613
	pesos_i(5517) := b"0000000000000000_0000000000000000_0101001000010110_0010100010000000"; -- 0.3206506073474884
	pesos_i(5518) := b"0000000000000000_0000000000000000_0100011001010100_0001100010000000"; -- 0.274720698595047
	pesos_i(5519) := b"1111111111111111_1111111111111111_1000110100000010_0101001110000000"; -- -0.44918325543403625
	pesos_i(5520) := b"1111111111111111_1111111111111111_1110110001011011_1100001110000000"; -- -0.07672479748725891
	pesos_i(5521) := b"0000000000000000_0000000000000000_0100000100111001_1001110010000000"; -- 0.25478532910346985
	pesos_i(5522) := b"0000000000000000_0000000000000000_0001011111101100_0110011100000000"; -- 0.09345096349716187
	pesos_i(5523) := b"0000000000000000_0000000000000000_0101111110000000_1111100100000000"; -- 0.3730617165565491
	pesos_i(5524) := b"0000000000000000_0000000000000000_0010110111101110_1001111110000000"; -- 0.17942234873771667
	pesos_i(5525) := b"0000000000000000_0000000000000000_0010000011011110_0010101001000000"; -- 0.12838996946811676
	pesos_i(5526) := b"1111111111111111_1111111111111111_0100010100110110_0001001000000000"; -- -0.729643702507019
	pesos_i(5527) := b"1111111111111111_1111111111111111_1101001001101001_0101011110000000"; -- -0.17808011174201965
	pesos_i(5528) := b"1111111111111111_1111111111111111_1011110010011011_1111011010000000"; -- -0.26324519515037537
	pesos_i(5529) := b"1111111111111111_1111111111111111_1110010000111010_1111011110100000"; -- -0.1084752306342125
	pesos_i(5530) := b"1111111111111111_1111111111111111_1100111100010010_1011101000000000"; -- -0.19112050533294678
	pesos_i(5531) := b"0000000000000000_0000000000000000_0101001011000000_0100001010000000"; -- 0.32324615120887756
	pesos_i(5532) := b"0000000000000000_0000000000000000_0001010001110101_0011111000100000"; -- 0.07991398125886917
	pesos_i(5533) := b"0000000000000000_0000000000000000_0011011110100101_1110001111000000"; -- 0.2173750251531601
	pesos_i(5534) := b"1111111111111111_1111111111111111_1101011111100110_0100010010000000"; -- -0.15664264559745789
	pesos_i(5535) := b"0000000000000000_0000000000000000_0010001010000100_1011010111000000"; -- 0.13483749330043793
	pesos_i(5536) := b"1111111111111111_1111111111111111_1110101110110000_0011100010000000"; -- -0.07934233546257019
	pesos_i(5537) := b"1111111111111111_1111111111111111_1111110001011000_1110101011010000"; -- -0.014268230646848679
	pesos_i(5538) := b"0000000000000000_0000000000000000_0000111011100011_1011100111110000"; -- 0.058162327855825424
	pesos_i(5539) := b"0000000000000000_0000000000000000_0001010011001101_1001101010000000"; -- 0.0812622606754303
	pesos_i(5540) := b"0000000000000000_0000000000000000_0011110100010111_0011000010000000"; -- 0.2386350929737091
	pesos_i(5541) := b"0000000000000000_0000000000000000_0011000010011010_0011101001000000"; -- 0.18985332548618317
	pesos_i(5542) := b"1111111111111111_1111111111111111_1010010011101110_1101001010000000"; -- -0.3557308614253998
	pesos_i(5543) := b"1111111111111111_1111111111111111_1001101001010101_1010110100000000"; -- -0.39713019132614136
	pesos_i(5544) := b"1111111111111111_1111111111111111_0111011000101100_0010111000000000"; -- -0.5383883714675903
	pesos_i(5545) := b"0000000000000000_0000000000000000_0101010100101000_0001001010000000"; -- 0.33264270424842834
	pesos_i(5546) := b"0000000000000000_0000000000000000_0101011101011011_1100111100000000"; -- 0.341244637966156
	pesos_i(5547) := b"0000000000000000_0000000000000000_0001000001010111_0100110011100000"; -- 0.06383209675550461
	pesos_i(5548) := b"1111111111111111_1111111111111111_1111000111001101_1001101011000000"; -- -0.05545647442340851
	pesos_i(5549) := b"0000000000000000_0000000000000000_0001000001111001_0111001101000000"; -- 0.06435318291187286
	pesos_i(5550) := b"1111111111111111_1111111111111111_1010100001011010_0000100110000000"; -- -0.34237614274024963
	pesos_i(5551) := b"1111111111111111_1111111111111111_1101110000111101_1011010110000000"; -- -0.13968339562416077
	pesos_i(5552) := b"0000000000000000_0000000000000000_0000110000100001_0101001001010000"; -- 0.047383446246385574
	pesos_i(5553) := b"0000000000000000_0000000000000000_0111100000100101_0111000010000000"; -- 0.46932128071784973
	pesos_i(5554) := b"1111111111111111_1111111111111111_1100001100010001_1101101100000000"; -- -0.2380087971687317
	pesos_i(5555) := b"0000000000000000_0000000000000000_0000110011101011_0000100101000000"; -- 0.05046136677265167
	pesos_i(5556) := b"1111111111111111_1111111111111111_1100000101001111_1111000110000000"; -- -0.24487391114234924
	pesos_i(5557) := b"1111111111111111_1111111111111111_1011000001010100_1101001110000000"; -- -0.31120565533638
	pesos_i(5558) := b"0000000000000000_0000000000000000_0010110110111011_1001111110000000"; -- 0.17864415049552917
	pesos_i(5559) := b"1111111111111111_1111111111111111_1010001000110001_1101000000000000"; -- -0.3664274215698242
	pesos_i(5560) := b"0000000000000000_0000000000000000_0001110011101100_1000001011100000"; -- 0.11298387497663498
	pesos_i(5561) := b"1111111111111111_1111111111111111_1100111011011111_1110011100000000"; -- -0.19189602136611938
	pesos_i(5562) := b"0000000000000000_0000000000000000_0000001010000010_1100111111001000"; -- 0.009808527305722237
	pesos_i(5563) := b"0000000000000000_0000000000000000_0011001110000000_1000101100000000"; -- 0.20118016004562378
	pesos_i(5564) := b"1111111111111111_1111111111111111_1101101000100001_1010111101000000"; -- -0.1479235142469406
	pesos_i(5565) := b"0000000000000000_0000000000000000_0011010010100000_1100010000000000"; -- 0.20557808876037598
	pesos_i(5566) := b"0000000000000000_0000000000000000_0000110111101101_1101100100010000"; -- 0.05441052094101906
	pesos_i(5567) := b"0000000000000000_0000000000000000_0100011001000010_0111010000000000"; -- 0.27445149421691895
	pesos_i(5568) := b"1111111111111111_1111111111111111_1111101001010000_1001111110010000"; -- -0.022207286208868027
	pesos_i(5569) := b"0000000000000000_0000000000000000_0110111011111010_1010011000000000"; -- 0.4335120916366577
	pesos_i(5570) := b"0000000000000000_0000000000000000_0010001111001110_0001111110000000"; -- 0.13986393809318542
	pesos_i(5571) := b"1111111111111111_1111111111111111_1100110111010101_1101111110000000"; -- -0.1959553062915802
	pesos_i(5572) := b"1111111111111111_1111111111111111_1010111100100110_1100011100000000"; -- -0.3158145546913147
	pesos_i(5573) := b"0000000000000000_0000000000000000_0011100001011110_1001011011000000"; -- 0.2201933115720749
	pesos_i(5574) := b"0000000000000000_0000000000000000_0010100011010010_0111001010000000"; -- 0.15946117043495178
	pesos_i(5575) := b"0000000000000000_0000000000000000_0001110000101110_0101111000100000"; -- 0.11008251458406448
	pesos_i(5576) := b"1111111111111111_1111111111111111_1110111111111101_1011001111100000"; -- -0.06253505498170853
	pesos_i(5577) := b"0000000000000000_0000000000000000_0001111001010011_1100110111000000"; -- 0.11846624314785004
	pesos_i(5578) := b"0000000000000000_0000000000000000_0000111100010001_0010111110010000"; -- 0.05885598435997963
	pesos_i(5579) := b"0000000000000000_0000000000000000_0100111000101000_0000001100000000"; -- 0.3052980303764343
	pesos_i(5580) := b"0000000000000000_0000000000000000_0010100010000100_0100001111000000"; -- 0.15826819837093353
	pesos_i(5581) := b"1111111111111111_1111111111111111_1011111110101001_1001011010000000"; -- -0.2513185441493988
	pesos_i(5582) := b"1111111111111111_1111111111111111_1011100011001110_1100100110000000"; -- -0.27809467911720276
	pesos_i(5583) := b"0000000000000000_0000000000000000_0000010100111001_0110111011101000"; -- 0.02040761150419712
	pesos_i(5584) := b"0000000000000000_0000000000000000_0001110110011100_0011100001000000"; -- 0.11566497385501862
	pesos_i(5585) := b"1111111111111111_1111111111111111_1011000111100000_0000010110000000"; -- -0.30517545342445374
	pesos_i(5586) := b"0000000000000000_0000000000000000_0101110101011110_1110000010000000"; -- 0.3647289574146271
	pesos_i(5587) := b"0000000000000000_0000000000000000_0101101100001111_0011110000000000"; -- 0.355701208114624
	pesos_i(5588) := b"1111111111111111_1111111111111111_1110000110000001_0011001000100000"; -- -0.11912237852811813
	pesos_i(5589) := b"1111111111111111_1111111111111111_1100001000011101_0110001101000000"; -- -0.24173907935619354
	pesos_i(5590) := b"1111111111111111_1111111111111111_1101001111110111_1000111010000000"; -- -0.172003835439682
	pesos_i(5591) := b"0000000000000000_0000000000000000_0000100011100011_0111100001000000"; -- 0.03472091257572174
	pesos_i(5592) := b"1111111111111111_1111111111111111_1000000001110010_1111101110000000"; -- -0.498245507478714
	pesos_i(5593) := b"1111111111111111_1111111111111111_1101110000110000_0101111101000000"; -- -0.13988690078258514
	pesos_i(5594) := b"1111111111111111_1111111111111111_1101111001001110_1110001011000000"; -- -0.13160879909992218
	pesos_i(5595) := b"0000000000000000_0000000000000000_0001000111110000_1010010011100000"; -- 0.07007818669080734
	pesos_i(5596) := b"0000000000000000_0000000000000000_0111100110010000_1101010000000000"; -- 0.4748661518096924
	pesos_i(5597) := b"1111111111111111_1111111111111111_1111110000011001_1001101101001100"; -- -0.015234273858368397
	pesos_i(5598) := b"0000000000000000_0000000000000000_0000100000011001_1010000110010000"; -- 0.031641099601984024
	pesos_i(5599) := b"0000000000000000_0000000000000000_0011100111001001_1111011010000000"; -- 0.22573795914649963
	pesos_i(5600) := b"0000000000000000_0000000000000000_0011001001010001_1010100100000000"; -- 0.19655853509902954
	pesos_i(5601) := b"0000000000000000_0000000000000000_0001010001110101_0010110100100000"; -- 0.07991296797990799
	pesos_i(5602) := b"1111111111111111_1111111111111111_1100001110111111_0011111111000000"; -- -0.23536302149295807
	pesos_i(5603) := b"1111111111111111_1111111111111111_0010010010110010_0100011000000000"; -- -0.8566547632217407
	pesos_i(5604) := b"1111111111111111_1111111111111111_1100011111110100_0111000010000000"; -- -0.21892639994621277
	pesos_i(5605) := b"1111111111111111_1111111111111111_1111100011011001_0110001100000000"; -- -0.027932941913604736
	pesos_i(5606) := b"0000000000000000_0000000000000000_0001001100110110_0100100100000000"; -- 0.0750470757484436
	pesos_i(5607) := b"0000000000000000_0000000000000000_1000101000100101_1011101100000000"; -- 0.5396382212638855
	pesos_i(5608) := b"1111111111111111_1111111111111111_1111100011000000_0001111011001000"; -- -0.028318477794528008
	pesos_i(5609) := b"0000000000000000_0000000000000000_0101101000001000_1000000010000000"; -- 0.35169222950935364
	pesos_i(5610) := b"1111111111111111_1111111111111110_1010000110101110_0101100000000000"; -- -1.3684334754943848
	pesos_i(5611) := b"0000000000000000_0000000000000000_0000111000110010_0000000111010000"; -- 0.055450547486543655
	pesos_i(5612) := b"1111111111111111_1111111111111111_1101011000011110_0110001010000000"; -- -0.16359886527061462
	pesos_i(5613) := b"1111111111111111_1111111111111111_1011110000111010_0110010100000000"; -- -0.2647339701652527
	pesos_i(5614) := b"0000000000000000_0000000000000000_0101101101001000_1101111010000000"; -- 0.3565806448459625
	pesos_i(5615) := b"0000000000000000_0000000000000000_0100110101011001_0101001110000000"; -- 0.30214425921440125
	pesos_i(5616) := b"0000000000000000_0000000000000000_0100010010110000_1100000010000000"; -- 0.26832202076911926
	pesos_i(5617) := b"0000000000000000_0000000000000000_0100111000011101_0100000110000000"; -- 0.3051339089870453
	pesos_i(5618) := b"1111111111111111_1111111111111111_1101110110100011_0100111101000000"; -- -0.13422684371471405
	pesos_i(5619) := b"1111111111111111_1111111111111111_1100001111000101_0100100000000000"; -- -0.23527097702026367
	pesos_i(5620) := b"0000000000000000_0000000000000000_0101010011100000_1100001100000000"; -- 0.3315545916557312
	pesos_i(5621) := b"1111111111111111_1111111111111111_1101101010111111_1101010101000000"; -- -0.14551036059856415
	pesos_i(5622) := b"0000000000000000_0000000000000000_0101111100001100_1101010100000000"; -- 0.37128955125808716
	pesos_i(5623) := b"1111111111111111_1111111111111111_1110111001000101_1110001100100000"; -- -0.06924610584974289
	pesos_i(5624) := b"0000000000000000_0000000000000000_0100111000110011_0001001110000000"; -- 0.3054668605327606
	pesos_i(5625) := b"1111111111111111_1111111111111111_1011101011001100_1011111100000000"; -- -0.2703133225440979
	pesos_i(5626) := b"0000000000000000_0000000000000000_0011111110010000_1001011000000000"; -- 0.2482999563217163
	pesos_i(5627) := b"1111111111111111_1111111111111111_1001011000000011_0110000010000000"; -- -0.4140109717845917
	pesos_i(5628) := b"0000000000000000_0000000000000000_0001000011010000_1001010100000000"; -- 0.06568270921707153
	pesos_i(5629) := b"1111111111111111_1111111111111111_1101111110001101_1001101010000000"; -- -0.1267455518245697
	pesos_i(5630) := b"1111111111111111_1111111111111111_0100110101000000_0101000100000000"; -- -0.6982373595237732
	pesos_i(5631) := b"1111111111111111_1111111111111111_1110000000100100_1010101110000000"; -- -0.12444046139717102
	pesos_i(5632) := b"0000000000000000_0000000000000000_0001100011010010_0010100111100000"; -- 0.09695684164762497
	pesos_i(5633) := b"0000000000000000_0000000000000000_0010011110011000_1000110001000000"; -- 0.15467144548892975
	pesos_i(5634) := b"0000000000000000_0000000000000000_0010110111001111_0001100000000000"; -- 0.1789412498474121
	pesos_i(5635) := b"1111111111111111_1111111111111111_1111001000101011_1101111111100000"; -- -0.05401802808046341
	pesos_i(5636) := b"1111111111111111_1111111111111111_1101100011000110_0110100000000000"; -- -0.15322256088256836
	pesos_i(5637) := b"0000000000000000_0000000000000000_0001110100100100_1000110001000000"; -- 0.11383892595767975
	pesos_i(5638) := b"0000000000000000_0000000000000000_0010111001100100_1101001001000000"; -- 0.18122591078281403
	pesos_i(5639) := b"0000000000000000_0000000000000000_0110011011000001_0111000110000000"; -- 0.4013892114162445
	pesos_i(5640) := b"1111111111111111_1111111111111111_1101110110110010_1111111100000000"; -- -0.13398748636245728
	pesos_i(5641) := b"1111111111111111_1111111111111111_1010010001010010_0011100010000000"; -- -0.3581204116344452
	pesos_i(5642) := b"0000000000000000_0000000000000000_0000100011101011_0101010111000000"; -- 0.03484092652797699
	pesos_i(5643) := b"0000000000000000_0000000000000000_0011000100111111_0011010101000000"; -- 0.1923707276582718
	pesos_i(5644) := b"1111111111111111_1111111111111111_1100100111110001_1011101010000000"; -- -0.2111552655696869
	pesos_i(5645) := b"0000000000000000_0000000000000000_0101100111100000_1100101000000000"; -- 0.35108625888824463
	pesos_i(5646) := b"0000000000000000_0000000000000000_0101101101100010_0010001000000000"; -- 0.35696613788604736
	pesos_i(5647) := b"0000000000000000_0000000000000000_0011000011100101_0100000001000000"; -- 0.19099809229373932
	pesos_i(5648) := b"1111111111111111_1111111111111111_1111001011010111_0000000000100000"; -- -0.0514068529009819
	pesos_i(5649) := b"0000000000000000_0000000000000000_0100001101100011_1011001010000000"; -- 0.2632400095462799
	pesos_i(5650) := b"1111111111111111_1111111111111111_1100001010010001_0110010111000000"; -- -0.2399689108133316
	pesos_i(5651) := b"1111111111111111_1111111111111111_1110100110011101_1100011111100000"; -- -0.08743620663881302
	pesos_i(5652) := b"1111111111111111_1111111111111111_1110100111111101_1101110101000000"; -- -0.08597008883953094
	pesos_i(5653) := b"0000000000000000_0000000000000000_0110011110100110_0110110000000000"; -- 0.40488314628601074
	pesos_i(5654) := b"1111111111111111_1111111111111111_1110101011100101_1100101101100000"; -- -0.0824311152100563
	pesos_i(5655) := b"0000000000000000_0000000000000000_0000111010110100_1011110111100000"; -- 0.05744539946317673
	pesos_i(5656) := b"0000000000000000_0000000000000000_0010001000101000_1110100000000000"; -- 0.1334366798400879
	pesos_i(5657) := b"0000000000000000_0000000000000000_0010010101110001_0100111110000000"; -- 0.14626023173332214
	pesos_i(5658) := b"0000000000000000_0000000000000000_0010011000110110_1111000011000000"; -- 0.14927582442760468
	pesos_i(5659) := b"1111111111111111_1111111111111111_1010011110001110_1011100000000000"; -- -0.34547853469848633
	pesos_i(5660) := b"1111111111111111_1111111111111111_1110010000101101_1000110011100000"; -- -0.10867995768785477
	pesos_i(5661) := b"1111111111111111_1111111111111111_1111000100001001_0011000101110000"; -- -0.05845347419381142
	pesos_i(5662) := b"1111111111111111_1111111111111111_1101101101000000_0010111100000000"; -- -0.14355188608169556
	pesos_i(5663) := b"1111111111111111_1111111111111111_1100001001000111_0011001001000000"; -- -0.24110113084316254
	pesos_i(5664) := b"0000000000000000_0000000000000000_0111101010101000_0101111110000000"; -- 0.47913166880607605
	pesos_i(5665) := b"0000000000000000_0000000000000000_0101010000111111_1101111000000000"; -- 0.32909953594207764
	pesos_i(5666) := b"1111111111111111_1111111111111111_1100001001010111_1011000000000000"; -- -0.24084949493408203
	pesos_i(5667) := b"1111111111111111_1111111111111111_1100100001001111_1100101110000000"; -- -0.2175324261188507
	pesos_i(5668) := b"0000000000000000_0000000000000000_0011111111101000_0110100001000000"; -- 0.24964000284671783
	pesos_i(5669) := b"0000000000000000_0000000000000000_0010111000000010_0111101110000000"; -- 0.17972537875175476
	pesos_i(5670) := b"1111111111111111_1111111111111111_1100111101110101_0101000001000000"; -- -0.18961618840694427
	pesos_i(5671) := b"0000000000000000_0000000000000000_0000110010001011_0110111001110000"; -- 0.04900255426764488
	pesos_i(5672) := b"1111111111111111_1111111111111111_1100110111010011_0000100100000000"; -- -0.19599860906600952
	pesos_i(5673) := b"1111111111111111_1111111111111111_1101100000011010_0110001001000000"; -- -0.15584741532802582
	pesos_i(5674) := b"0000000000000000_0000000000000000_0010001101000010_1111110111000000"; -- 0.13774095475673676
	pesos_i(5675) := b"0000000000000000_0000000000000000_0110110010001100_0011001100000000"; -- 0.42401427030563354
	pesos_i(5676) := b"1111111111111111_1111111111111111_1111011111011010_0100001101010000"; -- -0.031825821846723557
	pesos_i(5677) := b"1111111111111111_1111111111111111_1111111110010111_1000011010101001"; -- -0.0015941464807838202
	pesos_i(5678) := b"0000000000000000_0000000000000000_0001110000100011_0010110000100000"; -- 0.10991168767213821
	pesos_i(5679) := b"1111111111111111_1111111111111111_1011011011101000_1111101100000000"; -- -0.2855075001716614
	pesos_i(5680) := b"1111111111111111_1111111111111111_1111000011110011_0111011010000000"; -- -0.058785051107406616
	pesos_i(5681) := b"0000000000000000_0000000000000000_0100110100001010_1110101000000000"; -- 0.30094778537750244
	pesos_i(5682) := b"1111111111111111_1111111111111111_1111000111011110_1100001111100000"; -- -0.05519462376832962
	pesos_i(5683) := b"0000000000000000_0000000000000000_0100000101111100_0000110000000000"; -- 0.2557990550994873
	pesos_i(5684) := b"1111111111111111_1111111111111111_1101110010001010_0111011111000000"; -- -0.13851214945316315
	pesos_i(5685) := b"1111111111111111_1111111111111111_1110010100010110_0100110110100000"; -- -0.10512842983007431
	pesos_i(5686) := b"0000000000000000_0000000000000000_0001110001100110_1000111000000000"; -- 0.1109398603439331
	pesos_i(5687) := b"1111111111111111_1111111111111111_1110111000011101_1001000010000000"; -- -0.06986138224601746
	pesos_i(5688) := b"1111111111111111_1111111111111111_1110001001001000_0110011100100000"; -- -0.11608272045850754
	pesos_i(5689) := b"0000000000000000_0000000000000000_0000101001000101_1001101100100000"; -- 0.04012460261583328
	pesos_i(5690) := b"1111111111111111_1111111111111111_1111111011001011_0111110110001100"; -- -0.004707482643425465
	pesos_i(5691) := b"0000000000000000_0000000000000000_0001101111101011_1011100011100000"; -- 0.10906558483839035
	pesos_i(5692) := b"1111111111111111_1111111111111111_1111101110110011_0011111011110000"; -- -0.01679617539048195
	pesos_i(5693) := b"1111111111111111_1111111111111111_1101100100111111_1010011100000000"; -- -0.151372492313385
	pesos_i(5694) := b"0000000000000000_0000000000000000_0010010101001010_1000100100000000"; -- 0.14566856622695923
	pesos_i(5695) := b"0000000000000000_0000000000000000_0101111101110110_0100000110000000"; -- 0.3728981912136078
	pesos_i(5696) := b"0000000000000000_0000000000000000_0001010110010011_1100110010000000"; -- 0.08428648114204407
	pesos_i(5697) := b"0000000000000000_0000000000000000_0100000100001110_0011110010000000"; -- 0.2541234791278839
	pesos_i(5698) := b"0000000000000000_0000000000000000_0001010001000111_0011101000000000"; -- 0.07921183109283447
	pesos_i(5699) := b"1111111111111111_1111111111111111_1111000001010010_0001101101010000"; -- -0.06124715134501457
	pesos_i(5700) := b"0000000000000000_0000000000000000_0010100001000010_0101110010000000"; -- 0.15726259350776672
	pesos_i(5701) := b"0000000000000000_0000000000000000_0100011001000001_0100000010000000"; -- 0.2744331657886505
	pesos_i(5702) := b"0000000000000000_0000000000000000_0001001110000010_1101010111100000"; -- 0.07621514052152634
	pesos_i(5703) := b"1111111111111111_1111111111111111_1110101010111110_1101000111000000"; -- -0.08302582800388336
	pesos_i(5704) := b"0000000000000000_0000000000000000_0010101110100011_1100111110000000"; -- 0.1704683005809784
	pesos_i(5705) := b"1111111111111111_1111111111111111_1101101001001100_1101101001000000"; -- -0.14726482331752777
	pesos_i(5706) := b"0000000000000000_0000000000000000_0010110100100101_1001000111000000"; -- 0.1763545125722885
	pesos_i(5707) := b"0000000000000000_0000000000000000_0100010100000001_1101100010000000"; -- 0.26955941319465637
	pesos_i(5708) := b"1111111111111111_1111111111111111_1100010111010001_0101011000000000"; -- -0.22727453708648682
	pesos_i(5709) := b"1111111111111111_1111111111111111_1111101000111101_0011100111000000"; -- -0.02250327169895172
	pesos_i(5710) := b"0000000000000000_0000000000000000_1000101010111000_0100001100000000"; -- 0.5418741106987
	pesos_i(5711) := b"0000000000000000_0000000000000000_0101010110110000_0111000010000000"; -- 0.33472350239753723
	pesos_i(5712) := b"0000000000000000_0000000000000000_0100111100101101_0001001100000000"; -- 0.30928152799606323
	pesos_i(5713) := b"0000000000000000_0000000000000000_0001011110011001_1001001100100000"; -- 0.09218711405992508
	pesos_i(5714) := b"0000000000000000_0000000000000000_0011011001010011_0100101001000000"; -- 0.21220840513706207
	pesos_i(5715) := b"0000000000000000_0000000000000000_0001111110111001_1110110101100000"; -- 0.12393077462911606
	pesos_i(5716) := b"0000000000000000_0000000000000000_0001000101110101_1010110001100000"; -- 0.06820180267095566
	pesos_i(5717) := b"0000000000000000_0000000000000000_0001111000111010_1100000111000000"; -- 0.11808405816555023
	pesos_i(5718) := b"0000000000000000_0000000000000000_0110001000011000_1111011100000000"; -- 0.3831934332847595
	pesos_i(5719) := b"0000000000000000_0000000000000000_0100010100011101_0000110100000000"; -- 0.2699745297431946
	pesos_i(5720) := b"1111111111111111_1111111111111111_1100001000111001_1101011011000000"; -- -0.24130494892597198
	pesos_i(5721) := b"0000000000000000_0000000000000000_0001100100000111_0011011010100000"; -- 0.09776631742715836
	pesos_i(5722) := b"0000000000000000_0000000000000000_0000100001000100_1101110000010000"; -- 0.032300714403390884
	pesos_i(5723) := b"1111111111111111_1111111111111111_1111100111101011_0010111001101000"; -- -0.023755168542265892
	pesos_i(5724) := b"0000000000000000_0000000000000000_0000101110011101_1010011101110000"; -- 0.04537435993552208
	pesos_i(5725) := b"0000000000000000_0000000000000000_0001011101001001_0111110010100000"; -- 0.09096506983041763
	pesos_i(5726) := b"1111111111111111_1111111111111111_1101110101111111_0101101000000000"; -- -0.13477551937103271
	pesos_i(5727) := b"0000000000000000_0000000000000000_0100110000000010_0001111110000000"; -- 0.2969073951244354
	pesos_i(5728) := b"1111111111111111_1111111111111111_1111011000100011_1000110001000000"; -- -0.03852008283138275
	pesos_i(5729) := b"0000000000000000_0000000000000000_0000110100010111_0110000001010000"; -- 0.05113794282078743
	pesos_i(5730) := b"0000000000000000_0000000000000000_0010011011111001_0101101000000000"; -- 0.15224230289459229
	pesos_i(5731) := b"1111111111111111_1111111111111111_1101001000001110_1000101001000000"; -- -0.1794656366109848
	pesos_i(5732) := b"1111111111111111_1111111111111111_1100110101000100_0100011010000000"; -- -0.19817695021629333
	pesos_i(5733) := b"1111111111111111_1111111111111111_1100011111001111_0101010111000000"; -- -0.219492569565773
	pesos_i(5734) := b"0000000000000000_0000000000000000_0010010001111000_1000101110000000"; -- 0.14246436953544617
	pesos_i(5735) := b"1111111111111111_1111111111111111_1110011011011000_1010100001100000"; -- -0.09825656563043594
	pesos_i(5736) := b"0000000000000000_0000000000000000_0000011010100111_0111010101001000"; -- 0.025992708280682564
	pesos_i(5737) := b"1111111111111111_1111111111111111_1111001110110010_0011011011000000"; -- -0.04806192219257355
	pesos_i(5738) := b"0000000000000000_0000000000000000_0001110111011100_0110010110100000"; -- 0.1166442409157753
	pesos_i(5739) := b"0000000000000000_0000000000000000_0010011111110011_1111001100000000"; -- 0.15606611967086792
	pesos_i(5740) := b"0000000000000000_0000000000000000_0001100011011110_0110000010000000"; -- 0.09714320302009583
	pesos_i(5741) := b"0000000000000000_0000000000000000_0010110010001011_1111010011000000"; -- 0.17401055991649628
	pesos_i(5742) := b"1111111111111111_1111111111111111_1111001111001001_0000011101000000"; -- -0.04771380126476288
	pesos_i(5743) := b"0000000000000000_0000000000000000_0001010111101010_0010011111100000"; -- 0.08560418337583542
	pesos_i(5744) := b"0000000000000000_0000000000000000_0001101010100100_1100101010100000"; -- 0.10407701879739761
	pesos_i(5745) := b"1111111111111111_1111111111111111_1100100110100011_1000001010000000"; -- -0.2123487889766693
	pesos_i(5746) := b"0000000000000000_0000000000000000_0010110101011000_0101110011000000"; -- 0.17712955176830292
	pesos_i(5747) := b"0000000000000000_0000000000000000_0111000110000100_0010110100000000"; -- 0.4434230923652649
	pesos_i(5748) := b"1111111111111111_1111111111111111_1110001110101100_0001001011000000"; -- -0.11065562069416046
	pesos_i(5749) := b"0000000000000000_0000000000000000_0010100000010001_0111100010000000"; -- 0.15651658177375793
	pesos_i(5750) := b"0000000000000000_0000000000000000_0111001111110010_1110101000000000"; -- 0.45292532444000244
	pesos_i(5751) := b"0000000000000000_0000000000000000_0000100101110001_1000111000110000"; -- 0.0368889681994915
	pesos_i(5752) := b"0000000000000000_0000000000000000_0111010110000010_0101001110000000"; -- 0.45901986956596375
	pesos_i(5753) := b"0000000000000000_0000000000000000_0011100001011100_1011101111000000"; -- 0.22016499936580658
	pesos_i(5754) := b"0000000000000000_0000000000000000_0011001101100001_1100110101000000"; -- 0.20071108639240265
	pesos_i(5755) := b"0000000000000000_0000000000000000_0010100101010001_0010100110000000"; -- 0.16139468550682068
	pesos_i(5756) := b"0000000000000000_0000000000000000_0011000011001101_0001000101000000"; -- 0.19062907993793488
	pesos_i(5757) := b"0000000000000000_0000000000000000_0001010001011100_1011001110000000"; -- 0.07953950762748718
	pesos_i(5758) := b"1111111111111111_1111111111111111_1101100000100100_0000101100000000"; -- -0.15570002794265747
	pesos_i(5759) := b"0000000000000000_0000000000000000_0010111110101110_0001111110000000"; -- 0.18625065684318542
	pesos_i(5760) := b"0000000000000000_0000000000000000_0011000100111001_1000110000000000"; -- 0.19228434562683105
	pesos_i(5761) := b"0000000000000000_0000000000000000_0000011001011100_1111011010110000"; -- 0.02485601231455803
	pesos_i(5762) := b"0000000000000000_0000000000000000_0000100111010000_1011111001110000"; -- 0.03834142908453941
	pesos_i(5763) := b"0000000000000000_0000000000000000_0010011011111111_0111011010000000"; -- 0.15233555436134338
	pesos_i(5764) := b"1111111111111111_1111111111111111_1010100100000010_1001011100000000"; -- -0.3398042321205139
	pesos_i(5765) := b"1111111111111111_1111111111111111_1101110110011111_0001110111000000"; -- -0.13429082930088043
	pesos_i(5766) := b"0000000000000000_0000000000000000_0010011111101011_1101010100000000"; -- 0.15594226121902466
	pesos_i(5767) := b"1111111111111111_1111111111111111_1111010011100111_1010100011110000"; -- -0.04334015026688576
	pesos_i(5768) := b"1111111111111111_1111111111111111_0111010101001101_1000101000000000"; -- -0.5417855978012085
	pesos_i(5769) := b"1111111111111111_1111111111111111_1011111011110001_0011011000000000"; -- -0.25413191318511963
	pesos_i(5770) := b"0000000000000000_0000000000000000_0011111111001001_0000010010000000"; -- 0.249161034822464
	pesos_i(5771) := b"0000000000000000_0000000000000000_0010101001011010_0111001100000000"; -- 0.16544264554977417
	pesos_i(5772) := b"0000000000000000_0000000000000000_0001000111011100_1010101001000000"; -- 0.06977333128452301
	pesos_i(5773) := b"0000000000000000_0000000000000000_0100010011111010_1101110010000000"; -- 0.269452840089798
	pesos_i(5774) := b"0000000000000000_0000000000000000_0101011111001011_0000101100000000"; -- 0.34294193983078003
	pesos_i(5775) := b"0000000000000000_0000000000000000_0000011110001001_0001010111011000"; -- 0.029435506090521812
	pesos_i(5776) := b"1111111111111111_1111111111111111_1101111011000101_0100111100000000"; -- -0.12980180978775024
	pesos_i(5777) := b"0000000000000000_0000000000000000_0100101110010010_1011010010000000"; -- 0.29520729184150696
	pesos_i(5778) := b"1111111111111111_1111111111111111_1100001011011011_1111001001000000"; -- -0.23883138597011566
	pesos_i(5779) := b"0000000000000000_0000000000000000_0001001010011000_0000010111100000"; -- 0.07263218611478806
	pesos_i(5780) := b"0000000000000000_0000000000000000_0100010100101001_0010001010000000"; -- 0.27015891671180725
	pesos_i(5781) := b"0000000000000000_0000000000000000_0000100011000111_0110101101110000"; -- 0.034292902797460556
	pesos_i(5782) := b"0000000000000000_0000000000000000_0000101101001011_1110001001010000"; -- 0.04412664845585823
	pesos_i(5783) := b"0000000000000000_0000000000000000_0010000100010110_0010001100000000"; -- 0.12924402952194214
	pesos_i(5784) := b"1111111111111111_1111111111111111_1110010010110011_0100001010000000"; -- -0.10663971304893494
	pesos_i(5785) := b"1111111111111111_1111111111111111_1101111011001011_1001111010000000"; -- -0.1297055184841156
	pesos_i(5786) := b"0000000000000000_0000000000000000_0010010101100000_1111000010000000"; -- 0.14601042866706848
	pesos_i(5787) := b"1111111111111111_1111111111111111_1100010101000000_1100011101000000"; -- -0.2294803112745285
	pesos_i(5788) := b"0000000000000000_0000000000000000_0000010100101101_1000110001111000"; -- 0.020226268097758293
	pesos_i(5789) := b"1111111111111111_1111111111111111_1110010110111111_0001111110100000"; -- -0.10255243629217148
	pesos_i(5790) := b"1111111111111111_1111111111111111_1110111000001000_1000010010100000"; -- -0.07018252462148666
	pesos_i(5791) := b"1111111111111111_1111111111111111_1110000111110000_0010000011100000"; -- -0.11742968112230301
	pesos_i(5792) := b"1111111111111111_1111111111111111_1111100000001000_1000111111111000"; -- -0.031119348481297493
	pesos_i(5793) := b"0000000000000000_0000000000000000_0010010010101011_0100011010000000"; -- 0.14323845505714417
	pesos_i(5794) := b"0000000000000000_0000000000000000_0000110000111010_0001001101000000"; -- 0.047761157155036926
	pesos_i(5795) := b"1111111111111111_1111111111111111_1101110011001010_0001111100000000"; -- -0.13754087686538696
	pesos_i(5796) := b"1111111111111111_1111111111111111_1110100110010011_1101101000000000"; -- -0.08758771419525146
	pesos_i(5797) := b"0000000000000000_0000000000000000_0001110110100010_0101001010000000"; -- 0.11575809121131897
	pesos_i(5798) := b"0000000000000000_0000000000000000_0001000100100010_1100000010100000"; -- 0.06693653017282486
	pesos_i(5799) := b"1111111111111111_1111111111111111_1111100111000011_1011110111100000"; -- -0.024356968700885773
	pesos_i(5800) := b"0000000000000000_0000000000000000_0100100100011010_0010100000000000"; -- 0.285555362701416
	pesos_i(5801) := b"0000000000000000_0000000000000000_0100000010010001_1101100000000000"; -- 0.252225399017334
	pesos_i(5802) := b"0000000000000000_0000000000000000_0001101110111010_1110001101100000"; -- 0.1083204373717308
	pesos_i(5803) := b"1111111111111111_1111111111111111_1110110001100111_1010000111000000"; -- -0.07654370367527008
	pesos_i(5804) := b"1111111111111111_1111111111111111_1111100011010010_1010110100011000"; -- -0.02803533710539341
	pesos_i(5805) := b"0000000000000000_0000000000000000_0010000111100001_0110000000000000"; -- 0.13234519958496094
	pesos_i(5806) := b"1111111111111111_1111111111111111_1000111101010011_1111101100000000"; -- -0.4401248097419739
	pesos_i(5807) := b"0000000000000000_0000000000000000_0000111001110010_1000111010000000"; -- 0.05643549561500549
	pesos_i(5808) := b"0000000000000000_0000000000000000_0011110100000100_1101111010000000"; -- 0.23835554718971252
	pesos_i(5809) := b"1111111111111111_1111111111111111_1101111001001001_0101111010000000"; -- -0.13169297575950623
	pesos_i(5810) := b"1111111111111111_1111111111111111_1110100111010011_1111110000100000"; -- -0.0866091176867485
	pesos_i(5811) := b"0000000000000000_0000000000000000_0010010010011000_0011000101000000"; -- 0.1429472714662552
	pesos_i(5812) := b"0000000000000000_0000000000000000_0000110111011001_1001010100000000"; -- 0.05410128831863403
	pesos_i(5813) := b"1111111111111111_1111111111111111_1001001010001110_1001111110000000"; -- -0.4275112450122833
	pesos_i(5814) := b"0000000000000000_0000000000000000_0011001111110110_0100101011000000"; -- 0.20297686755657196
	pesos_i(5815) := b"0000000000000000_0000000000000000_0000001101111011_0010001100110000"; -- 0.013597678393125534
	pesos_i(5816) := b"1111111111111111_1111111111111111_1100110010110000_0100111011000000"; -- -0.20043475925922394
	pesos_i(5817) := b"0000000000000000_0000000000000000_0100111001111101_1011001100000000"; -- 0.3066055178642273
	pesos_i(5818) := b"0000000000000000_0000000000000000_0001110111000000_1000010111000000"; -- 0.11621890962123871
	pesos_i(5819) := b"0000000000000000_0000000000000000_0100111011100001_0011111000000000"; -- 0.3081244230270386
	pesos_i(5820) := b"1111111111111111_1111111111111111_1110111100100101_1101011000100000"; -- -0.06582891196012497
	pesos_i(5821) := b"1111111111111111_1111111111111111_1111101101000111_0010110010010000"; -- -0.018445219844579697
	pesos_i(5822) := b"0000000000000000_0000000000000000_0010111110101100_1110101101000000"; -- 0.1862322837114334
	pesos_i(5823) := b"0000000000000000_0000000000000000_0000010001100000_1000101111001000"; -- 0.01709817536175251
	pesos_i(5824) := b"0000000000000000_0000000000000000_0010111101000110_0000011100000000"; -- 0.18466228246688843
	pesos_i(5825) := b"1111111111111111_1111111111111111_1110100011000100_0111111001100000"; -- -0.09075174480676651
	pesos_i(5826) := b"1111111111111111_1111111111111111_1111101010010111_1000101110011000"; -- -0.021125102415680885
	pesos_i(5827) := b"0000000000000000_0000000000000000_0000011110100000_1100111011101000"; -- 0.029797488823533058
	pesos_i(5828) := b"1111111111111111_1111111111111111_1110101101001001_0010111110000000"; -- -0.08091452717781067
	pesos_i(5829) := b"0000000000000000_0000000000000000_0000100111100100_0111000101010000"; -- 0.03864200785756111
	pesos_i(5830) := b"1111111111111111_1111111111111111_0111001111101110_1001000000000000"; -- -0.5471410751342773
	pesos_i(5831) := b"1111111111111111_1111111111111111_1011000110110101_0101110000000000"; -- -0.30582642555236816
	pesos_i(5832) := b"0000000000000000_0000000000000000_0000100010001100_0110011110010000"; -- 0.03339240327477455
	pesos_i(5833) := b"1111111111111111_1111111111111111_1100010001111110_0010110100000000"; -- -0.2324497103691101
	pesos_i(5834) := b"1111111111111111_1111111111111111_1011110101010101_0011100010000000"; -- -0.2604183852672577
	pesos_i(5835) := b"0000000000000000_0000000000000000_0001000111100110_0111110000000000"; -- 0.06992316246032715
	pesos_i(5836) := b"1111111111111111_1111111111111111_1100010010000001_1011110100000000"; -- -0.23239535093307495
	pesos_i(5837) := b"0000000000000000_0000000000000000_0001101111011010_0001111000000000"; -- 0.10879695415496826
	pesos_i(5838) := b"0000000000000000_0000000000000000_0010001011100010_0000010011000000"; -- 0.13626126945018768
	pesos_i(5839) := b"1111111111111111_1111111111111111_1100010001010100_1001011010000000"; -- -0.2330842912197113
	pesos_i(5840) := b"1111111111111111_1111111111111111_1101010011000101_0001110110000000"; -- -0.16886726021766663
	pesos_i(5841) := b"1111111111111111_1111111111111111_1110111001010100_1100101010000000"; -- -0.06901869177818298
	pesos_i(5842) := b"0000000000000000_0000000000000000_0001010101111110_0011101010000000"; -- 0.08395734429359436
	pesos_i(5843) := b"0000000000000000_0000000000000000_0010011110000100_0100001100000000"; -- 0.15436190366744995
	pesos_i(5844) := b"1111111111111111_1111111111111111_1011100111100110_1000000010000000"; -- -0.27382656931877136
	pesos_i(5845) := b"1111111111111111_1111111111111111_1111011100000010_0001110001000000"; -- -0.035124048590660095
	pesos_i(5846) := b"0000000000000000_0000000000000000_0000011110100001_0000000111000000"; -- 0.029800519347190857
	pesos_i(5847) := b"1111111111111111_1111111111111111_1010000011010010_1011011000000000"; -- -0.3717848062515259
	pesos_i(5848) := b"0000000000000000_0000000000000000_0000101101001110_1001010011010000"; -- 0.04416780546307564
	pesos_i(5849) := b"0000000000000000_0000000000000000_0011010100000010_1000100111000000"; -- 0.2070699781179428
	pesos_i(5850) := b"1111111111111111_1111111111111111_1011000100100100_0100101000000000"; -- -0.3080400228500366
	pesos_i(5851) := b"1111111111111111_1111111111111111_1111001001101111_1010100110010000"; -- -0.05298366770148277
	pesos_i(5852) := b"1111111111111111_1111111111111111_1110111010110101_1111101000000000"; -- -0.06753575801849365
	pesos_i(5853) := b"1111111111111111_1111111111111111_1101110001110110_1111000101000000"; -- -0.13881008327007294
	pesos_i(5854) := b"0000000000000000_0000000000000000_0100000100000000_1011010110000000"; -- 0.25391706824302673
	pesos_i(5855) := b"0000000000000000_0000000000000000_0100110100011110_0010110110000000"; -- 0.3012417256832123
	pesos_i(5856) := b"1111111111111111_1111111111111111_1011010011100101_0111001000000000"; -- -0.2933739423751831
	pesos_i(5857) := b"1111111111111111_1111111111111111_1101101001001011_1111010001000000"; -- -0.1472785323858261
	pesos_i(5858) := b"1111111111111111_1111111111111111_1101101100110000_1111010110000000"; -- -0.14378419518470764
	pesos_i(5859) := b"0000000000000000_0000000000000000_0011011101000111_1101110100000000"; -- 0.21594029664993286
	pesos_i(5860) := b"0000000000000000_0000000000000000_0011010011110010_1000110000000000"; -- 0.20682597160339355
	pesos_i(5861) := b"0000000000000000_0000000000000000_0010111100011011_0011010101000000"; -- 0.1840089112520218
	pesos_i(5862) := b"0000000000000000_0000000000000000_0001100001011011_0101110111000000"; -- 0.09514413774013519
	pesos_i(5863) := b"0000000000000000_0000000000000000_0010010110101111_0111011001000000"; -- 0.1472085863351822
	pesos_i(5864) := b"1111111111111111_1111111111111111_1111000001001011_1100010000000000"; -- -0.06134390830993652
	pesos_i(5865) := b"1111111111111111_1111111111111111_1110010111101000_0110101110100000"; -- -0.10192229598760605
	pesos_i(5866) := b"0000000000000000_0000000000000000_0001110010111010_1011011111100000"; -- 0.11222409456968307
	pesos_i(5867) := b"1111111111111111_1111111111111111_1110011011110101_0110100011000000"; -- -0.09781785309314728
	pesos_i(5868) := b"0000000000000000_0000000000000000_0100101100100010_0100101000000000"; -- 0.2934919595718384
	pesos_i(5869) := b"0000000000000000_0000000000000000_0001011011101010_0101011010100000"; -- 0.08951321989297867
	pesos_i(5870) := b"1111111111111111_1111111111111111_1110100110101011_1010010110000000"; -- -0.08722463250160217
	pesos_i(5871) := b"0000000000000000_0000000000000000_0000010100001110_0010111111011000"; -- 0.019747724756598473
	pesos_i(5872) := b"1111111111111111_1111111111111111_1010110100110110_0100111000000000"; -- -0.3233901262283325
	pesos_i(5873) := b"1111111111111111_1111111111111111_1111100001100100_0101010011001000"; -- -0.029719067737460136
	pesos_i(5874) := b"0000000000000000_0000000000000000_0001110110011111_1011011110000000"; -- 0.11571833491325378
	pesos_i(5875) := b"1111111111111111_1111111111111111_1110111001010001_0101111010000000"; -- -0.06907090544700623
	pesos_i(5876) := b"1111111111111111_1111111111111111_1011100111010100_1001011100000000"; -- -0.2740998864173889
	pesos_i(5877) := b"0000000000000000_0000000000000000_0001101011111100_1001010011100000"; -- 0.10541658848524094
	pesos_i(5878) := b"0000000000000000_0000000000000000_0100010110011110_1010000100000000"; -- 0.27195173501968384
	pesos_i(5879) := b"0000000000000000_0000000000000000_0100101111100110_0011100100000000"; -- 0.2964816689491272
	pesos_i(5880) := b"0000000000000000_0000000000000000_0001100111010001_1110110110000000"; -- 0.10085949301719666
	pesos_i(5881) := b"0000000000000000_0000000000000000_0101000111100111_1001011110000000"; -- 0.31994006037712097
	pesos_i(5882) := b"1111111111111111_1111111111111111_1101111001000100_0111001100000000"; -- -0.13176804780960083
	pesos_i(5883) := b"0000000000000000_0000000000000000_0000001111000001_0110110000000000"; -- 0.014670133590698242
	pesos_i(5884) := b"0000000000000000_0000000000000000_0001011101010000_1001011001100000"; -- 0.0910734161734581
	pesos_i(5885) := b"1111111111111111_1111111111111111_1101101011001001_0111011101000000"; -- -0.14536337554454803
	pesos_i(5886) := b"0000000000000000_0000000000000000_0001110010110100_0000101001100000"; -- 0.11212220042943954
	pesos_i(5887) := b"1111111111111111_1111111111111111_1100100111100100_1111001011000000"; -- -0.21135027706623077
	pesos_i(5888) := b"0000000000000000_0000000000000000_0100010110101011_0001111110000000"; -- 0.2721423804759979
	pesos_i(5889) := b"1111111111111111_1111111111111111_1101110011001010_0010101001000000"; -- -0.13754020631313324
	pesos_i(5890) := b"1111111111111111_1111111111111111_1110101011110000_0000000011000000"; -- -0.08227534592151642
	pesos_i(5891) := b"1111111111111111_1111111111111111_1110100101011001_1001000000100000"; -- -0.08847712725400925
	pesos_i(5892) := b"1111111111111111_1111111111111111_1011010110101100_0001010100000000"; -- -0.2903429865837097
	pesos_i(5893) := b"1111111111111111_1111111111111111_1111011001100101_1011110011010000"; -- -0.03751010820269585
	pesos_i(5894) := b"0000000000000000_0000000000000000_0100111110111101_0110000010000000"; -- 0.3114834129810333
	pesos_i(5895) := b"1111111111111111_1111111111111111_1111010011000110_0101000011000000"; -- -0.04384894669055939
	pesos_i(5896) := b"1111111111111111_1111111111111111_0101100110000101_1000000100000000"; -- -0.6503066420555115
	pesos_i(5897) := b"0000000000000000_0000000000000000_0100010001001100_1010010000000000"; -- 0.26679444313049316
	pesos_i(5898) := b"0000000000000000_0000000000000000_0000010010101010_0001010010100000"; -- 0.018220223486423492
	pesos_i(5899) := b"1111111111111111_1111111111111111_1101101100111111_1000000011000000"; -- -0.14356227219104767
	pesos_i(5900) := b"0000000000000000_0000000000000000_0001010111001011_0101011100100000"; -- 0.08513397723436356
	pesos_i(5901) := b"0000000000000000_0000000000000000_0000000010100101_0111011001011011"; -- 0.0025247547309845686
	pesos_i(5902) := b"0000000000000000_0000000000000000_0001101000110000_1100110000100000"; -- 0.10230708867311478
	pesos_i(5903) := b"1111111111111111_1111111111111111_1111110001101010_1011011000000000"; -- -0.013996720314025879
	pesos_i(5904) := b"0000000000000000_0000000000000000_0001111110010001_0110100000000000"; -- 0.12331247329711914
	pesos_i(5905) := b"0000000000000000_0000000000000000_0010010010100100_1010000010000000"; -- 0.14313700795173645
	pesos_i(5906) := b"1111111111111111_1111111111111111_1111110110011000_1000111001101100"; -- -0.00939092505723238
	pesos_i(5907) := b"0000000000000000_0000000000000000_0101100001100010_0111001000000000"; -- 0.3452521562576294
	pesos_i(5908) := b"0000000000000000_0000000000000000_0001011110010100_1010101111000000"; -- 0.09211228787899017
	pesos_i(5909) := b"0000000000000000_0000000000000000_0000110101000110_0001001111010000"; -- 0.05185054615139961
	pesos_i(5910) := b"0000000000000000_0000000000000000_0001011011000000_1100011111000000"; -- 0.08887909352779388
	pesos_i(5911) := b"1111111111111111_1111111111111111_1101110111111110_1010101101000000"; -- -0.13283281028270721
	pesos_i(5912) := b"1111111111111111_1111111111111111_1100010010011100_1010101001000000"; -- -0.231984481215477
	pesos_i(5913) := b"0000000000000000_0000000000000000_0001011000110100_0101101101100000"; -- 0.08673640340566635
	pesos_i(5914) := b"0000000000000000_0000000000000000_0011110000111110_0010001110000000"; -- 0.23532316088676453
	pesos_i(5915) := b"1111111111111111_1111111111111111_1111010110000111_1010110111110000"; -- -0.04089844599366188
	pesos_i(5916) := b"1111111111111111_1111111111111111_1101100100011101_0011100100000000"; -- -0.1518978476524353
	pesos_i(5917) := b"1111111111111111_1111111111111111_1110011010010110_1111011101000000"; -- -0.09925894439220428
	pesos_i(5918) := b"0000000000000000_0000000000000000_0000110100000011_0010001101000000"; -- 0.05082912743091583
	pesos_i(5919) := b"1111111111111111_1111111111111111_1101010001011011_1000001110000000"; -- -0.17047861218452454
	pesos_i(5920) := b"1111111111111111_1111111111111111_1110011000001100_1101010110000000"; -- -0.10136666893959045
	pesos_i(5921) := b"0000000000000000_0000000000000000_0001110111010101_0001011001100000"; -- 0.11653270572423935
	pesos_i(5922) := b"0000000000000000_0000000000000000_0000000111110011_0100000111010100"; -- 0.007618059404194355
	pesos_i(5923) := b"1111111111111111_1111111111111111_1111100000010100_0001110011111000"; -- -0.030943097546696663
	pesos_i(5924) := b"1111111111111111_1111111111111111_1100111001100100_1101101101000000"; -- -0.193773552775383
	pesos_i(5925) := b"0000000000000000_0000000000000000_0110001101111001_0011010010000000"; -- 0.3885681927204132
	pesos_i(5926) := b"1111111111111111_1111111111111111_1110101110000111_1101000011000000"; -- -0.07995887100696564
	pesos_i(5927) := b"0000000000000000_0000000000000000_0001001011111101_1111111001000000"; -- 0.07418812811374664
	pesos_i(5928) := b"0000000000000000_0000000000000000_0010010000100111_1101010010000000"; -- 0.14123275876045227
	pesos_i(5929) := b"0000000000000000_0000000000000000_0001011100000111_0110111001000000"; -- 0.08995713293552399
	pesos_i(5930) := b"0000000000000000_0000000000000000_0000010111010101_0111100010000000"; -- 0.022788554430007935
	pesos_i(5931) := b"1111111111111111_1111111111111111_1101110101110000_1010000101000000"; -- -0.13500015437602997
	pesos_i(5932) := b"0000000000000000_0000000000000000_0000010011100010_1001000110110000"; -- 0.019082169979810715
	pesos_i(5933) := b"1111111111111111_1111111111111111_1111111010011100_0010110110111110"; -- -0.005429402459412813
	pesos_i(5934) := b"1111111111111111_1111111111111111_1001000110001101_1101001010000000"; -- -0.4314297139644623
	pesos_i(5935) := b"0000000000000000_0000000000000000_0001110110010101_1010011010000000"; -- 0.1155647337436676
	pesos_i(5936) := b"0000000000000000_0000000000000000_0011000010000101_1101000101000000"; -- 0.18954189121723175
	pesos_i(5937) := b"0000000000000000_0000000000000000_0001010000000111_1000001010000000"; -- 0.07823958992958069
	pesos_i(5938) := b"1111111111111111_1111111111111111_1110101101111101_1101000000100000"; -- -0.08011149615049362
	pesos_i(5939) := b"1111111111111111_1111111111111111_1111010101100100_0010000001010000"; -- -0.041440945118665695
	pesos_i(5940) := b"1111111111111111_1111111111111111_1111010101000000_1101000100100000"; -- -0.041979722678661346
	pesos_i(5941) := b"1111111111111111_1111111111111111_1101000000110001_1100010010000000"; -- -0.18674060702323914
	pesos_i(5942) := b"0000000000000000_0000000000000000_0000011011010010_1100011010110000"; -- 0.02665368840098381
	pesos_i(5943) := b"0000000000000000_0000000000000000_0001001111010001_0100110111100000"; -- 0.07741247862577438
	pesos_i(5944) := b"0000000000000000_0000000000000000_0000001011100001_1110110000100000"; -- 0.011259801685810089
	pesos_i(5945) := b"0000000000000000_0000000000000000_0001001101101010_0001000110100000"; -- 0.07583723217248917
	pesos_i(5946) := b"1111111111111111_1111111111111111_1111011010001000_0001101100010000"; -- -0.036985691636800766
	pesos_i(5947) := b"0000000000000000_0000000000000000_0000101110101110_0101000111010000"; -- 0.04562865570187569
	pesos_i(5948) := b"0000000000000000_0000000000000000_0001110111011000_0101100110000000"; -- 0.1165824830532074
	pesos_i(5949) := b"0000000000000000_0000000000000000_0010100001101011_0011101100000000"; -- 0.15788620710372925
	pesos_i(5950) := b"1111111111111111_1111111111111111_1111001100101111_0010000000000000"; -- -0.05006217956542969
	pesos_i(5951) := b"0000000000000000_0000000000000000_0010000011001010_0000111101000000"; -- 0.12808318436145782
	pesos_i(5952) := b"0000000000000000_0000000000000000_0001100001010001_1101111001000000"; -- 0.09499920904636383
	pesos_i(5953) := b"1111111111111111_1111111111111111_1110001110011101_0111110100000000"; -- -0.11087816953659058
	pesos_i(5954) := b"0000000000000000_0000000000000000_0100000010000011_0100011000000000"; -- 0.2520030736923218
	pesos_i(5955) := b"0000000000000000_0000000000000000_0001010111011011_1001101110100000"; -- 0.08538220077753067
	pesos_i(5956) := b"1111111111111111_1111111111111111_1110010100000110_0111000011000000"; -- -0.10537047684192657
	pesos_i(5957) := b"1111111111111111_1111111111111111_1111010011111000_0100111101100000"; -- -0.04308608919382095
	pesos_i(5958) := b"1111111111111111_1111111111111111_1000011001101011_1101101000000000"; -- -0.47491681575775146
	pesos_i(5959) := b"1111111111111111_1111111111111111_1111000000001000_1100111100010000"; -- -0.062365587800741196
	pesos_i(5960) := b"1111111111111111_1111111111111111_1111111000000011_1110100101100010"; -- -0.007752812933176756
	pesos_i(5961) := b"1111111111111111_1111111111111111_1111001111111101_0100111000010000"; -- -0.04691612347960472
	pesos_i(5962) := b"1111111111111111_1111111111111111_1110001010001000_1011100000000000"; -- -0.11510133743286133
	pesos_i(5963) := b"0000000000000000_0000000000000000_0011011000010100_1101011000000000"; -- 0.21125543117523193
	pesos_i(5964) := b"0000000000000000_0000000000000000_0011001110001001_0000001101000000"; -- 0.20130939781665802
	pesos_i(5965) := b"0000000000000000_0000000000000000_0000010100110011_0101111001110000"; -- 0.020315077155828476
	pesos_i(5966) := b"0000000000000000_0000000000000000_0001100010001010_0100110000100000"; -- 0.09586025029420853
	pesos_i(5967) := b"1111111111111111_1111111111111111_1011110000100110_1100011110000000"; -- -0.2650332748889923
	pesos_i(5968) := b"0000000000000000_0000000000000000_0001100000101101_1111001100000000"; -- 0.09445112943649292
	pesos_i(5969) := b"1111111111111111_1111111111111111_1111111111101010_1011111011101001"; -- -0.0003243141691200435
	pesos_i(5970) := b"0000000000000000_0000000000000000_0010010111011101_1111010011000000"; -- 0.14791803061962128
	pesos_i(5971) := b"0000000000000000_0000000000000000_0000111101110110_1110010011010000"; -- 0.06040792539715767
	pesos_i(5972) := b"1111111111111111_1111111111111111_1100001111010001_1101100100000000"; -- -0.23507922887802124
	pesos_i(5973) := b"1111111111111111_1111111111111111_1111000010110001_0100100011100000"; -- -0.05979485064744949
	pesos_i(5974) := b"1111111111111111_1111111111111111_1110010110001101_1001001111100000"; -- -0.10330844670534134
	pesos_i(5975) := b"1111111111111111_1111111111111111_1101111010010010_0110001000000000"; -- -0.130578875541687
	pesos_i(5976) := b"1111111111111111_1111111111111111_1111010100100111_0000110000100000"; -- -0.0423729345202446
	pesos_i(5977) := b"0000000000000000_0000000000000000_0001001101110111_1101010100000000"; -- 0.07604724168777466
	pesos_i(5978) := b"0000000000000000_0000000000000000_0000001100111100_0111111111000100"; -- 0.01264189276844263
	pesos_i(5979) := b"0000000000000000_0000000000000000_0011000100001110_0001000000000000"; -- 0.1916208267211914
	pesos_i(5980) := b"0000000000000000_0000000000000000_0101110010100000_1010111010000000"; -- 0.3618268072605133
	pesos_i(5981) := b"0000000000000000_0000000000000000_0011000110010101_0011100001000000"; -- 0.19368316233158112
	pesos_i(5982) := b"1111111111111111_1111111111111111_1110011111001010_0110010111100000"; -- -0.09456790238618851
	pesos_i(5983) := b"0000000000000000_0000000000000000_0000110000001110_1110001111100000"; -- 0.04710220545530319
	pesos_i(5984) := b"0000000000000000_0000000000000000_0000110110100101_0111011000110000"; -- 0.05330599471926689
	pesos_i(5985) := b"1111111111111111_1111111111111111_1111010011111001_0000010000110000"; -- -0.0430753119289875
	pesos_i(5986) := b"1111111111111111_1111111111111111_0101010101001111_1111000100000000"; -- -0.6667489409446716
	pesos_i(5987) := b"0000000000000000_0000000000000000_0001110000010010_0010011000100000"; -- 0.10965193063020706
	pesos_i(5988) := b"0000000000000000_0000000000000000_0000101010100001_0001000011010000"; -- 0.041520167142152786
	pesos_i(5989) := b"1111111111111111_1111111111111111_1111110001001001_1110100010000100"; -- -0.014497249387204647
	pesos_i(5990) := b"1111111111111111_1111111111111111_1110101101010010_0000010011000000"; -- -0.08077974617481232
	pesos_i(5991) := b"0000000000000000_0000000000000000_0011011101100110_0111101010000000"; -- 0.21640744805335999
	pesos_i(5992) := b"0000000000000000_0000000000000000_0010110011110000_0011111000000000"; -- 0.17554080486297607
	pesos_i(5993) := b"1111111111111111_1111111111111111_1100000110111111_1001011000000000"; -- -0.2431703805923462
	pesos_i(5994) := b"0000000000000000_0000000000000000_0000000100010011_1111001111011010"; -- 0.0042107016779482365
	pesos_i(5995) := b"0000000000000000_0000000000000000_0010001110011001_1111100101000000"; -- 0.13906820118427277
	pesos_i(5996) := b"0000000000000000_0000000000000000_0000101101110001_1001011110010000"; -- 0.04470202699303627
	pesos_i(5997) := b"1111111111111111_1111111111111111_1011001111111101_1101000100000000"; -- -0.29690831899642944
	pesos_i(5998) := b"0000000000000000_0000000000000000_0010110100101101_1011101101000000"; -- 0.1764790564775467
	pesos_i(5999) := b"1111111111111111_1111111111111111_1110101011001110_1001100100100000"; -- -0.08278506249189377
	pesos_i(6000) := b"1111111111111111_1111111111111111_1011101100110001_1010000000000000"; -- -0.26877403259277344
	pesos_i(6001) := b"0000000000000000_0000000000000000_0101010010100011_0001111000000000"; -- 0.33061397075653076
	pesos_i(6002) := b"0000000000000000_0000000000000000_0010011100011010_1100101100000000"; -- 0.1527525782585144
	pesos_i(6003) := b"1111111111111111_1111111111111111_1100111111001000_1111100100000000"; -- -0.18833965063095093
	pesos_i(6004) := b"0000000000000000_0000000000000000_0001001101100111_0100001100000000"; -- 0.07579439878463745
	pesos_i(6005) := b"1111111111111111_1111111111111111_1101000010000000_0000010001000000"; -- -0.1855466216802597
	pesos_i(6006) := b"0000000000000000_0000000000000000_0000101100010000_1000111101010000"; -- 0.04322143271565437
	pesos_i(6007) := b"0000000000000000_0000000000000000_0010010110100010_1100111111000000"; -- 0.1470155566930771
	pesos_i(6008) := b"1111111111111111_1111111111111111_1111111101010101_0001100010100011"; -- -0.002607784466817975
	pesos_i(6009) := b"1111111111111111_1111111111111111_1111110010100110_0001101000010100"; -- -0.013090486638247967
	pesos_i(6010) := b"1111111111111111_1111111111111111_1101100001101100_1010010110000000"; -- -0.15459218621253967
	pesos_i(6011) := b"1111111111111111_1111111111111111_1111001100010100_1001011101000000"; -- -0.05046705901622772
	pesos_i(6012) := b"0000000000000000_0000000000000000_0011101010000111_0101011110000000"; -- 0.22862765192985535
	pesos_i(6013) := b"1111111111111111_1111111111111111_1101000010101011_0110110110000000"; -- -0.1848842203617096
	pesos_i(6014) := b"0000000000000000_0000000000000000_0000011010110111_0000110100111000"; -- 0.026230646297335625
	pesos_i(6015) := b"1111111111111111_1111111111111111_1110010001110001_1101000100100000"; -- -0.10763829201459885
	pesos_i(6016) := b"0000000000000000_0000000000000000_0011001110011000_0011010011000000"; -- 0.2015412300825119
	pesos_i(6017) := b"1111111111111111_1111111111111111_1110000111100111_0010011011000000"; -- -0.11756666004657745
	pesos_i(6018) := b"0000000000000000_0000000000000000_0000001011110110_0011101110100100"; -- 0.011569716967642307
	pesos_i(6019) := b"0000000000000000_0000000000000000_0000111000000001_1101101110110000"; -- 0.054715853184461594
	pesos_i(6020) := b"0000000000000000_0000000000000000_0000101011001110_1011111110010000"; -- 0.042217228561639786
	pesos_i(6021) := b"0000000000000000_0000000000000000_0001110011011100_0101111000100000"; -- 0.11273754388093948
	pesos_i(6022) := b"0000000000000000_0000000000000000_0000101100000110_1110010010110000"; -- 0.04307393357157707
	pesos_i(6023) := b"0000000000000000_0000000000000000_0010010111010110_1110111000000000"; -- 0.14781081676483154
	pesos_i(6024) := b"1111111111111111_1111111111111111_1100100000011110_0100000011000000"; -- -0.2182883769273758
	pesos_i(6025) := b"0000000000000000_0000000000000000_0000011110000010_0101101011110000"; -- 0.029332812875509262
	pesos_i(6026) := b"1111111111111111_1111111111111111_1011111011000000_0011110100000000"; -- -0.2548791766166687
	pesos_i(6027) := b"1111111111111111_1111111111111111_1100101000111001_1110000110000000"; -- -0.21005430817604065
	pesos_i(6028) := b"1111111111111111_1111111111111111_1110010100110010_0011010100100000"; -- -0.10470264405012131
	pesos_i(6029) := b"0000000000000000_0000000000000000_0010101000010110_0010010110000000"; -- 0.16440042853355408
	pesos_i(6030) := b"1111111111111111_1111111111111111_1011110010000111_1100011000000000"; -- -0.263553261756897
	pesos_i(6031) := b"0000000000000000_0000000000000000_0000001010011111_1010101000010000"; -- 0.010248783975839615
	pesos_i(6032) := b"0000000000000000_0000000000000000_0000000111110011_0111111100001000"; -- 0.007621707394719124
	pesos_i(6033) := b"1111111111111111_1111111111111111_1111000101010111_1000001100010000"; -- -0.057258423417806625
	pesos_i(6034) := b"0000000000000000_0000000000000000_0001001100010110_0101111110000000"; -- 0.07456013560295105
	pesos_i(6035) := b"0000000000000000_0000000000000000_0000101010000010_0100010111110000"; -- 0.04105031117796898
	pesos_i(6036) := b"0000000000000000_0000000000000000_0001111001000110_1011101100100000"; -- 0.1182667687535286
	pesos_i(6037) := b"1111111111111111_1111111111111111_1110011100011110_0110001100000000"; -- -0.09719258546829224
	pesos_i(6038) := b"0000000000000000_0000000000000000_0000010101011110_1111111111001000"; -- 0.020980821922421455
	pesos_i(6039) := b"0000000000000000_0000000000000000_0000000011100111_0111011000111110"; -- 0.0035318280570209026
	pesos_i(6040) := b"1111111111111111_1111111111111111_1101100011010010_0001101111000000"; -- -0.15304400026798248
	pesos_i(6041) := b"1111111111111111_1111111111111111_1110011100001011_1111101010000000"; -- -0.09747347235679626
	pesos_i(6042) := b"0000000000000000_0000000000000000_0000101111010100_0101100011110000"; -- 0.04620891436934471
	pesos_i(6043) := b"0000000000000000_0000000000000000_0001110100010110_1110111111000000"; -- 0.1136312335729599
	pesos_i(6044) := b"0000000000000000_0000000000000000_0010000011010010_0101110101000000"; -- 0.1282099038362503
	pesos_i(6045) := b"0000000000000000_0000000000000000_0010101111001010_0100110111000000"; -- 0.1710556596517563
	pesos_i(6046) := b"1111111111111111_1111111111111111_1110111011001111_0111110001000000"; -- -0.06714652478694916
	pesos_i(6047) := b"0000000000000000_0000000000000000_0001010010110000_0001111110100000"; -- 0.08081243187189102
	pesos_i(6048) := b"0000000000000000_0000000000000000_0000011100011010_0011101010100000"; -- 0.027743972837924957
	pesos_i(6049) := b"0000000000000000_0000000000000000_0001110001001010_1001010001000000"; -- 0.11051298677921295
	pesos_i(6050) := b"0000000000000000_0000000000000000_0000001110010110_0001110100010100"; -- 0.01400930155068636
	pesos_i(6051) := b"1111111111111111_1111111111111111_1110110101110011_0101011011100000"; -- -0.07245881110429764
	pesos_i(6052) := b"0000000000000000_0000000000000000_0000000100001001_0001001100111000"; -- 0.004044724628329277
	pesos_i(6053) := b"1111111111111111_1111111111111111_1110110111100111_1000110100000000"; -- -0.07068556547164917
	pesos_i(6054) := b"1111111111111111_1111111111111111_1101010000100111_0110000011000000"; -- -0.17127414047718048
	pesos_i(6055) := b"0000000000000000_0000000000000000_0001101000101001_1100101011000000"; -- 0.10220019519329071
	pesos_i(6056) := b"0000000000000000_0000000000000000_0000110111111001_0001101001100000"; -- 0.05458226054906845
	pesos_i(6057) := b"0000000000000000_0000000000000000_0010011001010011_1001100001000000"; -- 0.14971305429935455
	pesos_i(6058) := b"1111111111111111_1111111111111111_1111100000000110_0011010011100000"; -- -0.0311552956700325
	pesos_i(6059) := b"1111111111111111_1111111111111111_1110110001010010_1001100001000000"; -- -0.07686470448970795
	pesos_i(6060) := b"0000000000000000_0000000000000000_0001111111000011_1000011000000000"; -- 0.1240772008895874
	pesos_i(6061) := b"1111111111111111_1111111111111111_1101100000100000_1110111101000000"; -- -0.1557474583387375
	pesos_i(6062) := b"1111111111111111_1111111111111111_1100101011110100_1110011100000000"; -- -0.20720058679580688
	pesos_i(6063) := b"0000000000000000_0000000000000000_0010001000001000_1101000001000000"; -- 0.13294698297977448
	pesos_i(6064) := b"1111111111111111_1111111111111111_1101011000011101_0001100101000000"; -- -0.16361849009990692
	pesos_i(6065) := b"0000000000000000_0000000000000000_0010100010001111_0010000001000000"; -- 0.1584339290857315
	pesos_i(6066) := b"1111111111111111_1111111111111111_1010100101100000_1111111010000000"; -- -0.33836373686790466
	pesos_i(6067) := b"0000000000000000_0000000000000000_0000111011011001_1010101001010000"; -- 0.05800880864262581
	pesos_i(6068) := b"1111111111111111_1111111111111111_1111011110010101_1111001010100000"; -- -0.03286822885274887
	pesos_i(6069) := b"0000000000000000_0000000000000000_0001001101100110_0001000011100000"; -- 0.07577615231275558
	pesos_i(6070) := b"1111111111111111_1111111111111111_1110111001110010_1001111100100000"; -- -0.06856351345777512
	pesos_i(6071) := b"0000000000000000_0000000000000000_0001010111001010_1001010111100000"; -- 0.08512245863676071
	pesos_i(6072) := b"1111111111111111_1111111111111111_1101010010111000_1010010100000000"; -- -0.16905754804611206
	pesos_i(6073) := b"0000000000000000_0000000000000000_0010010001000100_1011001010000000"; -- 0.1416732370853424
	pesos_i(6074) := b"1111111111111111_1111111111111111_1111101010011011_0001110110110000"; -- -0.02107061818242073
	pesos_i(6075) := b"1111111111111111_1111111111111111_1111010110000101_1100110000100000"; -- -0.04092716425657272
	pesos_i(6076) := b"0000000000000000_0000000000000000_0001001001100100_0011000110000000"; -- 0.07184132933616638
	pesos_i(6077) := b"0000000000000000_0000000000000000_0011101111011100_0101110000000000"; -- 0.23383116722106934
	pesos_i(6078) := b"0000000000000000_0000000000000000_0010010010111111_0110111001000000"; -- 0.143546000123024
	pesos_i(6079) := b"0000000000000000_0000000000000000_0001101100001111_1101001101000000"; -- 0.1057102233171463
	pesos_i(6080) := b"0000000000000000_0000000000000000_0011010111110111_0010100100000000"; -- 0.2108026146888733
	pesos_i(6081) := b"1111111111111111_1111111111111111_1100110011100011_0111100111000000"; -- -0.1996539980173111
	pesos_i(6082) := b"0000000000000000_0000000000000000_0011011110010010_1111100001000000"; -- 0.2170863300561905
	pesos_i(6083) := b"0000000000000000_0000000000000000_0010001010010010_1101100011000000"; -- 0.13505320250988007
	pesos_i(6084) := b"1111111111111111_1111111111111111_1010000101000100_0011111100000000"; -- -0.37005239725112915
	pesos_i(6085) := b"0000000000000000_0000000000000000_0001100101000111_0001101100100000"; -- 0.09874124079942703
	pesos_i(6086) := b"0000000000000000_0000000000000000_0010010111010110_0111001010000000"; -- 0.14780345559120178
	pesos_i(6087) := b"1111111111111111_1111111111111111_1110101111001011_0100000000000000"; -- -0.07892990112304688
	pesos_i(6088) := b"1111111111111111_1111111111111111_1110101001110011_1110111001000000"; -- -0.08416853845119476
	pesos_i(6089) := b"0000000000000000_0000000000000000_0000000100011110_0101001001010100"; -- 0.004368920810520649
	pesos_i(6090) := b"1111111111111111_1111111111111111_1010110100010101_0010101100000000"; -- -0.32389575242996216
	pesos_i(6091) := b"0000000000000000_0000000000000000_0000110100110010_0011110111010000"; -- 0.05154787376523018
	pesos_i(6092) := b"0000000000000000_0000000000000000_0010111011110110_0110111010000000"; -- 0.18344774842262268
	pesos_i(6093) := b"1111111111111111_1111111111111111_1110001000111011_0101100010000000"; -- -0.11628195643424988
	pesos_i(6094) := b"0000000000000000_0000000000000000_0010010000110111_0111000000000000"; -- 0.14147090911865234
	pesos_i(6095) := b"1111111111111111_1111111111111111_1111001111010011_0001000010100000"; -- -0.04756065458059311
	pesos_i(6096) := b"0000000000000000_0000000000000000_0001010000111111_1011110111000000"; -- 0.07909761369228363
	pesos_i(6097) := b"0000000000000000_0000000000000000_0011101011101001_1110110001000000"; -- 0.23013187944889069
	pesos_i(6098) := b"1111111111111111_1111111111111111_1111100011001100_0010010001101000"; -- -0.028135037049651146
	pesos_i(6099) := b"0000000000000000_0000000000000000_0011101110001000_1001110100000000"; -- 0.23255330324172974
	pesos_i(6100) := b"0000000000000000_0000000000000000_0001011100111010_0111110010100000"; -- 0.09073618799448013
	pesos_i(6101) := b"1111111111111111_1111111111111111_1101001001000110_0110001111000000"; -- -0.17861343920230865
	pesos_i(6102) := b"0000000000000000_0000000000000000_0000110001111001_1110010010110000"; -- 0.04873494431376457
	pesos_i(6103) := b"1111111111111111_1111111111111111_1011111110010010_1001001110000000"; -- -0.25166967511177063
	pesos_i(6104) := b"1111111111111111_1111111111111111_1111100100001000_1111011000010000"; -- -0.027207013219594955
	pesos_i(6105) := b"1111111111111111_1111111111111111_1110101010001110_0000001011100000"; -- -0.08377058058977127
	pesos_i(6106) := b"1111111111111111_1111111111111111_1110010100001101_0010111011100000"; -- -0.10526759177446365
	pesos_i(6107) := b"0000000000000000_0000000000000000_0011010010001100_0011010011000000"; -- 0.2052643746137619
	pesos_i(6108) := b"0000000000000000_0000000000000000_0010011000010110_1011100000000000"; -- 0.14878416061401367
	pesos_i(6109) := b"0000000000000000_0000000000000000_0010011011100011_1011011000000000"; -- 0.15191209316253662
	pesos_i(6110) := b"1111111111111111_1111111111111111_1111100010111000_0111110001001000"; -- -0.02843497507274151
	pesos_i(6111) := b"0000000000000000_0000000000000000_0000100110101001_0001100010110000"; -- 0.03773645684123039
	pesos_i(6112) := b"0000000000000000_0000000000000000_0001001111010001_1001101001000000"; -- 0.0774170309305191
	pesos_i(6113) := b"0000000000000000_0000000000000000_0010001001110110_0001011011000000"; -- 0.13461439311504364
	pesos_i(6114) := b"1111111111111111_1111111111111111_1100010011110100_1111011010000000"; -- -0.23063716292381287
	pesos_i(6115) := b"1111111111111111_1111111111111111_1011100011010111_0100101100000000"; -- -0.27796489000320435
	pesos_i(6116) := b"1111111111111111_1111111111111111_1110010000101101_0101111111100000"; -- -0.10868263989686966
	pesos_i(6117) := b"1111111111111111_1111111111111111_1100100000110010_0010001001000000"; -- -0.21798501908779144
	pesos_i(6118) := b"1111111111111111_1111111111111111_1101100101001010_0001001111000000"; -- -0.15121342241764069
	pesos_i(6119) := b"0000000000000000_0000000000000000_0010010000110101_0000101111000000"; -- 0.1414344161748886
	pesos_i(6120) := b"0000000000000000_0000000000000000_0000001101100010_0011000110011100"; -- 0.013217068277299404
	pesos_i(6121) := b"1111111111111111_1111111111111111_1100111111010000_1010111100000000"; -- -0.1882219910621643
	pesos_i(6122) := b"1111111111111111_1111111111111111_1111101110111111_0111101000110000"; -- -0.016609538346529007
	pesos_i(6123) := b"0000000000000000_0000000000000000_0010000111101011_1100001100000000"; -- 0.1325036883354187
	pesos_i(6124) := b"1111111111111111_1111111111111111_1111001000001100_0010001000010000"; -- -0.05450236424803734
	pesos_i(6125) := b"0000000000000000_0000000000000000_0000010110001000_0001101101111000"; -- 0.021608082577586174
	pesos_i(6126) := b"0000000000000000_0000000000000000_0010101010100111_0110100011000000"; -- 0.16661696135997772
	pesos_i(6127) := b"0000000000000000_0000000000000000_0000000011000101_1010100010010111"; -- 0.0030160301830619574
	pesos_i(6128) := b"0000000000000000_0000000000000000_0001110001001111_1010101011000000"; -- 0.1105906218290329
	pesos_i(6129) := b"0000000000000000_0000000000000000_0100001110100111_1111000010000000"; -- 0.264281302690506
	pesos_i(6130) := b"0000000000000000_0000000000000000_0011010000111110_1001000110000000"; -- 0.20407971739768982
	pesos_i(6131) := b"1111111111111111_1111111111111111_1100111110000001_0101011000000000"; -- -0.18943274021148682
	pesos_i(6132) := b"1111111111111111_1111111111111111_1111100110101000_0111010001110000"; -- -0.024773333221673965
	pesos_i(6133) := b"1111111111111111_1111111111111111_1111101011101010_1010001000100000"; -- -0.01985727995634079
	pesos_i(6134) := b"0000000000000000_0000000000000000_0001000010111000_1110100010100000"; -- 0.06532148271799088
	pesos_i(6135) := b"0000000000000000_0000000000000000_0000101001100011_0110111111000000"; -- 0.04057978093624115
	pesos_i(6136) := b"1111111111111111_1111111111111111_1110011001000110_0101010100100000"; -- -0.1004893109202385
	pesos_i(6137) := b"1111111111111111_1111111111111111_1101111111000100_0001011010000000"; -- -0.12591418623924255
	pesos_i(6138) := b"1111111111111111_1111111111111111_1101010011110101_0000001110000000"; -- -0.1681363880634308
	pesos_i(6139) := b"1111111111111111_1111111111111111_1010011110010110_1000101010000000"; -- -0.3453591763973236
	pesos_i(6140) := b"1111111111111111_1111111111111111_1111111110101010_1011000111010100"; -- -0.0013016563607379794
	pesos_i(6141) := b"1111111111111111_1111111111111111_1111001001010011_1101100111110000"; -- -0.05340803042054176
	pesos_i(6142) := b"0000000000000000_0000000000000000_0010101010110101_0111011011000000"; -- 0.16683141887187958
	pesos_i(6143) := b"1111111111111111_1111111111111111_1110011001111101_0010111000000000"; -- -0.09965240955352783
	pesos_i(6144) := b"0000000000000000_0000000000000000_0010111100100010_1100010010000000"; -- 0.18412426114082336
	pesos_i(6145) := b"0000000000000000_0000000000000000_0001101011001000_1100111010000000"; -- 0.10462656617164612
	pesos_i(6146) := b"0000000000000000_0000000000000000_0010101000011110_1110101101000000"; -- 0.1645342856645584
	pesos_i(6147) := b"1111111111111111_1111111111111111_1100101011010000_1110100000000000"; -- -0.2077498435974121
	pesos_i(6148) := b"0000000000000000_0000000000000000_0010110101111010_0010010000000000"; -- 0.17764496803283691
	pesos_i(6149) := b"1111111111111111_1111111111111111_1111000101001111_0111110101100000"; -- -0.057380832731723785
	pesos_i(6150) := b"0000000000000000_0000000000000000_0000101101010110_1100111111010000"; -- 0.044293392449617386
	pesos_i(6151) := b"1111111111111111_1111111111111111_1111111111100111_1101100010111001"; -- -0.0003685519623104483
	pesos_i(6152) := b"1111111111111111_1111111111111111_1110010001101111_0011101000100000"; -- -0.10767780989408493
	pesos_i(6153) := b"0000000000000000_0000000000000000_0000101001101000_1011011101010000"; -- 0.04066034033894539
	pesos_i(6154) := b"1111111111111111_1111111111111111_1111001010011100_0101101001100000"; -- -0.052301742136478424
	pesos_i(6155) := b"0000000000000000_0000000000000000_0000111111110111_1111000110000000"; -- 0.06237706542015076
	pesos_i(6156) := b"0000000000000000_0000000000000000_0000001010101011_1010100001001100"; -- 0.010431784205138683
	pesos_i(6157) := b"1111111111111111_1111111111111111_1111101100110001_1101011010110000"; -- -0.018770772963762283
	pesos_i(6158) := b"1111111111111111_1111111111111111_1110001101010101_1101000100000000"; -- -0.11197179555892944
	pesos_i(6159) := b"0000000000000000_0000000000000000_0001101100000011_0101001111000000"; -- 0.10551951825618744
	pesos_i(6160) := b"1111111111111111_1111111111111111_1100010110011010_0110110111000000"; -- -0.2281123548746109
	pesos_i(6161) := b"0000000000000000_0000000000000000_0100100100110111_0001101110000000"; -- 0.2859971225261688
	pesos_i(6162) := b"0000000000000000_0000000000000000_0010010100110000_0011100001000000"; -- 0.14526702463626862
	pesos_i(6163) := b"1111111111111111_1111111111111111_1101100000000001_1100010001000000"; -- -0.15622304379940033
	pesos_i(6164) := b"0000000000000000_0000000000000000_0010101110100011_0110001101000000"; -- 0.17046184837818146
	pesos_i(6165) := b"1111111111111111_1111111111111111_1111111011110101_1011011001010010"; -- -0.004063229542225599
	pesos_i(6166) := b"1111111111111111_1111111111111111_1111000001100110_0101110111010000"; -- -0.06093801185488701
	pesos_i(6167) := b"0000000000000000_0000000000000000_0010110010011110_0111100100000000"; -- 0.17429310083389282
	pesos_i(6168) := b"1111111111111111_1111111111111111_1111111010010101_1010011101101000"; -- -0.00552896223962307
	pesos_i(6169) := b"1111111111111111_1111111111111111_1111000100110100_0100010000110000"; -- -0.05779622867703438
	pesos_i(6170) := b"0000000000000000_0000000000000000_0100001101001010_1000100110000000"; -- 0.2628560960292816
	pesos_i(6171) := b"1111111111111111_1111111111111111_1101100110000000_0111011001000000"; -- -0.1503835767507553
	pesos_i(6172) := b"1111111111111111_1111111111111111_1111001010111111_0101100110010000"; -- -0.051767732948064804
	pesos_i(6173) := b"1111111111111111_1111111111111111_1101000000110101_1011000111000000"; -- -0.18668068945407867
	pesos_i(6174) := b"0000000000000000_0000000000000000_0010011000000000_0001011010000000"; -- 0.14843884110450745
	pesos_i(6175) := b"1111111111111111_1111111111111111_1110010011000011_0100100110100000"; -- -0.10639514774084091
	pesos_i(6176) := b"1111111111111111_1111111111111111_1111100100101011_0000001110101000"; -- -0.02668740414083004
	pesos_i(6177) := b"0000000000000000_0000000000000000_0011010010011101_0110000010000000"; -- 0.20552638173103333
	pesos_i(6178) := b"0000000000000000_0000000000000000_0001100001010001_0111111111000000"; -- 0.09499357640743256
	pesos_i(6179) := b"1111111111111111_1111111111111111_1110001010011010_1011011000000000"; -- -0.11482679843902588
	pesos_i(6180) := b"1111111111111111_1111111111111111_1111110100111101_1111000100100000"; -- -0.010773591697216034
	pesos_i(6181) := b"0000000000000000_0000000000000000_0010010101110000_1010001110000000"; -- 0.14624997973442078
	pesos_i(6182) := b"1111111111111111_1111111111111111_1100001111011111_0011100001000000"; -- -0.23487518727779388
	pesos_i(6183) := b"1111111111111111_1111111111111111_1111110000111110_0000010011000000"; -- -0.014678671956062317
	pesos_i(6184) := b"0000000000000000_0000000000000000_0001000011000100_1001100001000000"; -- 0.06549979746341705
	pesos_i(6185) := b"1111111111111111_1111111111111111_1101010111110101_1101001001000000"; -- -0.16421781480312347
	pesos_i(6186) := b"1111111111111111_1111111111111111_1100111000001011_1101000000000000"; -- -0.19513225555419922
	pesos_i(6187) := b"0000000000000000_0000000000000000_0000100100011001_1000100111000000"; -- 0.03554593026638031
	pesos_i(6188) := b"1111111111111111_1111111111111111_1101101110100101_0010011101000000"; -- -0.14201121032238007
	pesos_i(6189) := b"1111111111111111_1111111111111111_1111101100110101_0110110101111000"; -- -0.018716009333729744
	pesos_i(6190) := b"1111111111111111_1111111111111111_1011100110110100_1111000110000000"; -- -0.27458277344703674
	pesos_i(6191) := b"1111111111111111_1111111111111111_1101000011100111_0100011001000000"; -- -0.18397103250026703
	pesos_i(6192) := b"1111111111111111_1111111111111111_1110110111011010_1101110010100000"; -- -0.07087918370962143
	pesos_i(6193) := b"1111111111111111_1111111111111111_1101001000111001_0101000111000000"; -- -0.1788128763437271
	pesos_i(6194) := b"1111111111111111_1111111111111111_1111101000101101_1010101101001000"; -- -0.022740645334124565
	pesos_i(6195) := b"0000000000000000_0000000000000000_0000110110000111_1101000101100000"; -- 0.05285366624593735
	pesos_i(6196) := b"1111111111111111_1111111111111111_1101011111000101_1100000100000000"; -- -0.15713876485824585
	pesos_i(6197) := b"1111111111111111_1111111111111111_1101100010100100_0111101110000000"; -- -0.15374019742012024
	pesos_i(6198) := b"0000000000000000_0000000000000000_0010001010010101_1010100111000000"; -- 0.13509617745876312
	pesos_i(6199) := b"0000000000000000_0000000000000000_0000101111010111_0000111110110000"; -- 0.046250324696302414
	pesos_i(6200) := b"1111111111111111_1111111111111111_1101111110011010_1111000000000000"; -- -0.1265420913696289
	pesos_i(6201) := b"0000000000000000_0000000000000000_0011110110101000_0101000101000000"; -- 0.240849569439888
	pesos_i(6202) := b"1111111111111111_1111111111111111_1100100100011100_1101111100000000"; -- -0.2144032120704651
	pesos_i(6203) := b"0000000000000000_0000000000000000_0000111100011100_1010011101000000"; -- 0.059030964970588684
	pesos_i(6204) := b"0000000000000000_0000000000000000_0011010111001111_0111111110000000"; -- 0.21019741892814636
	pesos_i(6205) := b"0000000000000000_0000000000000000_0010010110011010_1001110100000000"; -- 0.14689046144485474
	pesos_i(6206) := b"0000000000000000_0000000000000000_0010000000011001_1010100111000000"; -- 0.12539158761501312
	pesos_i(6207) := b"0000000000000000_0000000000000000_0010000001001000_1010100011000000"; -- 0.12610869109630585
	pesos_i(6208) := b"0000000000000000_0000000000000000_0000110100111111_0100111100010000"; -- 0.051747266203165054
	pesos_i(6209) := b"0000000000000000_0000000000000000_0010101110011001_1000011001000000"; -- 0.1703113466501236
	pesos_i(6210) := b"1111111111111111_1111111111111111_1110011101110011_0101101011100000"; -- -0.09589607268571854
	pesos_i(6211) := b"0000000000000000_0000000000000000_0001111011010000_0110010011100000"; -- 0.12036734074354172
	pesos_i(6212) := b"0000000000000000_0000000000000000_0010000101111101_1100111001000000"; -- 0.13082589209079742
	pesos_i(6213) := b"1111111111111111_1111111111111111_1110100111000100_0011100100000000"; -- -0.0868496298789978
	pesos_i(6214) := b"1111111111111111_1111111111111111_1111101011110001_1101110010011000"; -- -0.01974698342382908
	pesos_i(6215) := b"1111111111111111_1111111111111111_1111110111000001_1101011011110000"; -- -0.00876099243760109
	pesos_i(6216) := b"0000000000000000_0000000000000000_0000001010000110_1010111011111100"; -- 0.009867607615888119
	pesos_i(6217) := b"1111111111111111_1111111111111111_1111010001011100_1110111001100000"; -- -0.045456983149051666
	pesos_i(6218) := b"1111111111111111_1111111111111111_1111010000111011_1010101101010000"; -- -0.045964520424604416
	pesos_i(6219) := b"0000000000000000_0000000000000000_0010001010010001_0010101000000000"; -- 0.13502752780914307
	pesos_i(6220) := b"0000000000000000_0000000000000000_0000001100011110_1000111001011000"; -- 0.012184998020529747
	pesos_i(6221) := b"1111111111111111_1111111111111111_1110110010111000_1000111010000000"; -- -0.0753088891506195
	pesos_i(6222) := b"0000000000000000_0000000000000000_0000110111001111_0100001110110000"; -- 0.053943853825330734
	pesos_i(6223) := b"1111111111111111_1111111111111111_1110001101100010_1101011111100000"; -- -0.11177302151918411
	pesos_i(6224) := b"1111111111111111_1111111111111111_1011101101000110_0000011000000000"; -- -0.26846277713775635
	pesos_i(6225) := b"0000000000000000_0000000000000000_0010111011110001_0111011010000000"; -- 0.18337193131446838
	pesos_i(6226) := b"1111111111111111_1111111111111111_1011101100000101_0001011010000000"; -- -0.26945361495018005
	pesos_i(6227) := b"0000000000000000_0000000000000000_0000101101010101_0100110000000000"; -- 0.04427027702331543
	pesos_i(6228) := b"0000000000000000_0000000000000000_0001010101100000_0100111000100000"; -- 0.08350075036287308
	pesos_i(6229) := b"0000000000000000_0000000000000000_0000111110010000_0010010100110000"; -- 0.060793232172727585
	pesos_i(6230) := b"0000000000000000_0000000000000000_0001111101000010_0000110100000000"; -- 0.12210160493850708
	pesos_i(6231) := b"1111111111111111_1111111111111111_1111110101011011_1110100100011000"; -- -0.010316306725144386
	pesos_i(6232) := b"0000000000000000_0000000000000000_0000000100011000_0011011111100100"; -- 0.0042757922783494
	pesos_i(6233) := b"0000000000000000_0000000000000000_0010101011001010_0010111000000000"; -- 0.16714751720428467
	pesos_i(6234) := b"0000000000000000_0000000000000000_0001010110100000_1110011011100000"; -- 0.08448641747236252
	pesos_i(6235) := b"1111111111111111_1111111111111111_1111000100111010_1111000010110000"; -- -0.05769439414143562
	pesos_i(6236) := b"1111111111111111_1111111111111111_1100010111000110_0101111110000000"; -- -0.22744181752204895
	pesos_i(6237) := b"1111111111111111_1111111111111111_1111110110010101_1011111000101000"; -- -0.00943385623395443
	pesos_i(6238) := b"1111111111111111_1111111111111111_1110010001001100_1101101011100000"; -- -0.10820228606462479
	pesos_i(6239) := b"0000000000000000_0000000000000000_0000011001011000_1100101110100000"; -- 0.02479241043329239
	pesos_i(6240) := b"1111111111111111_1111111111111111_1101111111000001_1111110111000000"; -- -0.12594617903232574
	pesos_i(6241) := b"0000000000000000_0000000000000000_0001100000001010_1101011001100000"; -- 0.09391536563634872
	pesos_i(6242) := b"1111111111111111_1111111111111111_1111010101100001_0010110010100000"; -- -0.0414859876036644
	pesos_i(6243) := b"0000000000000000_0000000000000000_0010011100110000_0011110110000000"; -- 0.1530798375606537
	pesos_i(6244) := b"0000000000000000_0000000000000000_0010110010111001_1101010010000000"; -- 0.17471054196357727
	pesos_i(6245) := b"0000000000000000_0000000000000000_0010001110010101_0001100010000000"; -- 0.1389937698841095
	pesos_i(6246) := b"1111111111111111_1111111111111111_1011000101010101_0000111010000000"; -- -0.30729588866233826
	pesos_i(6247) := b"0000000000000000_0000000000000000_0010101010010110_1101110000000000"; -- 0.16636443138122559
	pesos_i(6248) := b"1111111111111111_1111111111111111_1100100100011110_1011101010000000"; -- -0.2143748700618744
	pesos_i(6249) := b"0000000000000000_0000000000000000_0000100000110111_1110001001010000"; -- 0.03210272267460823
	pesos_i(6250) := b"0000000000000000_0000000000000000_0110011101001101_0100001010000000"; -- 0.40352264046669006
	pesos_i(6251) := b"0000000000000000_0000000000000000_0010101000100010_0001010010000000"; -- 0.1645825207233429
	pesos_i(6252) := b"1111111111111111_1111111111111111_1110001001111000_1011001101000000"; -- -0.11534576117992401
	pesos_i(6253) := b"0000000000000000_0000000000000000_0010010111101101_0110111100000000"; -- 0.14815419912338257
	pesos_i(6254) := b"1111111111111111_1111111111111111_1110101111011101_0000011110100000"; -- -0.07865860313177109
	pesos_i(6255) := b"1111111111111111_1111111111111111_1011100010110100_0100110100000000"; -- -0.2784988284111023
	pesos_i(6256) := b"1111111111111111_1111111111111111_1101101111111101_1000110000000000"; -- -0.14066243171691895
	pesos_i(6257) := b"0000000000000000_0000000000000000_0010001100111110_0001001111000000"; -- 0.13766597211360931
	pesos_i(6258) := b"0000000000000000_0000000000000000_0000101110011010_1100101101100000"; -- 0.045330725610256195
	pesos_i(6259) := b"0000000000000000_0000000000000000_0000110111010000_0000011101010000"; -- 0.05395551398396492
	pesos_i(6260) := b"1111111111111111_1111111111111111_1010000011111000_1110100000000000"; -- -0.3712019920349121
	pesos_i(6261) := b"0000000000000000_0000000000000000_0001010011100100_1001111001100000"; -- 0.0816134437918663
	pesos_i(6262) := b"1111111111111111_1111111111111111_1101111000000001_0010010110000000"; -- -0.13279500603675842
	pesos_i(6263) := b"0000000000000000_0000000000000000_0100001010100010_0011001100000000"; -- 0.26028746366500854
	pesos_i(6264) := b"1111111111111111_1111111111111111_1111000000110110_0010000001000000"; -- -0.061674103140830994
	pesos_i(6265) := b"0000000000000000_0000000000000000_0010010101110011_1111100000000000"; -- 0.1463007926940918
	pesos_i(6266) := b"1111111111111111_1111111111111111_1111100001100000_0110010100001000"; -- -0.029779134318232536
	pesos_i(6267) := b"0000000000000000_0000000000000000_0100000000110010_0000000110000000"; -- 0.25076302886009216
	pesos_i(6268) := b"0000000000000000_0000000000000000_0000001100101100_1001101001110000"; -- 0.0123993419110775
	pesos_i(6269) := b"1111111111111111_1111111111111111_1111000110001111_0011110101110000"; -- -0.05640808120369911
	pesos_i(6270) := b"0000000000000000_0000000000000000_0100010101101110_1110110110000000"; -- 0.27122387290000916
	pesos_i(6271) := b"0000000000000000_0000000000000000_0000010110110100_0001010101001000"; -- 0.022279100492596626
	pesos_i(6272) := b"1111111111111111_1111111111111111_1111000001001100_0101101010100000"; -- -0.06133493036031723
	pesos_i(6273) := b"1111111111111111_1111111111111111_1111111011011000_0001011111110100"; -- -0.0045151738449931145
	pesos_i(6274) := b"0000000000000000_0000000000000000_0011001101001111_1111110100000000"; -- 0.20043927431106567
	pesos_i(6275) := b"1111111111111111_1111111111111111_1101100010001010_1111010111000000"; -- -0.15412963926792145
	pesos_i(6276) := b"0000000000000000_0000000000000000_0011101000000010_0100110101000000"; -- 0.2265976220369339
	pesos_i(6277) := b"1111111111111111_1111111111111111_1101010101101100_0100101001000000"; -- -0.16631637513637543
	pesos_i(6278) := b"1111111111111111_1111111111111111_1101011101110111_0001000010000000"; -- -0.1583394706249237
	pesos_i(6279) := b"1111111111111111_1111111111111111_1010010110110111_1011110010000000"; -- -0.35266515612602234
	pesos_i(6280) := b"1111111111111111_1111111111111111_1111000101101100_1101100100110000"; -- -0.056932855397462845
	pesos_i(6281) := b"0000000000000000_0000000000000000_0001101010010101_0011011010000000"; -- 0.10383930802345276
	pesos_i(6282) := b"1111111111111111_1111111111111111_1011101101010110_0100111100000000"; -- -0.26821428537368774
	pesos_i(6283) := b"1111111111111111_1111111111111111_1110011110111111_0011010011000000"; -- -0.0947386771440506
	pesos_i(6284) := b"1111111111111111_1111111111111111_1110011011100001_0101101011000000"; -- -0.09812386333942413
	pesos_i(6285) := b"0000000000000000_0000000000000000_0000111101101000_0011111111100000"; -- 0.06018447130918503
	pesos_i(6286) := b"1111111111111111_1111111111111111_1111001011011101_0001011010110000"; -- -0.05131395533680916
	pesos_i(6287) := b"0000000000000000_0000000000000000_0000110000001001_1011011011000000"; -- 0.0470232218503952
	pesos_i(6288) := b"1111111111111111_1111111111111111_1011101101010000_0001001100000000"; -- -0.26830941438674927
	pesos_i(6289) := b"0000000000000000_0000000000000000_0011000011010010_0111100100000000"; -- 0.19071155786514282
	pesos_i(6290) := b"0000000000000000_0000000000000000_0000111011011111_1001000101100000"; -- 0.05809887498617172
	pesos_i(6291) := b"0000000000000000_0000000000000000_0010110101100100_0111111101000000"; -- 0.17731471359729767
	pesos_i(6292) := b"0000000000000000_0000000000000000_0000000100010111_0100101100111100"; -- 0.0042616864666342735
	pesos_i(6293) := b"0000000000000000_0000000000000000_0010000110111000_0111101101000000"; -- 0.13172121345996857
	pesos_i(6294) := b"0000000000000000_0000000000000000_0010101001110111_1110101001000000"; -- 0.16589225828647614
	pesos_i(6295) := b"0000000000000000_0000000000000000_0001000011100110_0111001000000000"; -- 0.0660163164138794
	pesos_i(6296) := b"1111111111111111_1111111111111111_1111000111001101_0100000110110000"; -- -0.055461782962083817
	pesos_i(6297) := b"1111111111111111_1111111111111111_1111101001110000_0111100011000000"; -- -0.02172131836414337
	pesos_i(6298) := b"0000000000000000_0000000000000000_0101001010001100_0111011100000000"; -- 0.32245582342147827
	pesos_i(6299) := b"0000000000000000_0000000000000000_0011001000110111_1101010000000000"; -- 0.19616436958312988
	pesos_i(6300) := b"1111111111111111_1111111111111111_1111100000100011_0100010001010000"; -- -0.03071187064051628
	pesos_i(6301) := b"0000000000000000_0000000000000000_0000000000000101_0001111110001100"; -- 7.817427103873342e-05
	pesos_i(6302) := b"0000000000000000_0000000000000000_0011110100111111_0101101101000000"; -- 0.23924799263477325
	pesos_i(6303) := b"1111111111111111_1111111111111111_1111100010000001_0010001110111000"; -- -0.02927948720753193
	pesos_i(6304) := b"0000000000000000_0000000000000000_0100100100100010_1110000110000000"; -- 0.28568848967552185
	pesos_i(6305) := b"1111111111111111_1111111111111111_1111101010110110_0011100110010000"; -- -0.020656969398260117
	pesos_i(6306) := b"0000000000000000_0000000000000000_0010111101110110_1110101011000000"; -- 0.18540827929973602
	pesos_i(6307) := b"0000000000000000_0000000000000000_0010000011110111_0000011001000000"; -- 0.12876929342746735
	pesos_i(6308) := b"1111111111111111_1111111111111111_1110110001000111_0010111000000000"; -- -0.07703888416290283
	pesos_i(6309) := b"0000000000000000_0000000000000000_0010101001101111_0100110111000000"; -- 0.1657608598470688
	pesos_i(6310) := b"1111111111111111_1111111111111111_1100110101001111_0011000110000000"; -- -0.19801035523414612
	pesos_i(6311) := b"1111111111111111_1111111111111111_1101010010010111_0110010000000000"; -- -0.16956496238708496
	pesos_i(6312) := b"0000000000000000_0000000000000000_0011111000110100_1010001110000000"; -- 0.24299070239067078
	pesos_i(6313) := b"1111111111111111_1111111111111111_1101111010111010_0100110101000000"; -- -0.1299697607755661
	pesos_i(6314) := b"1111111111111111_1111111111111111_1010111110010000_0111010110000000"; -- -0.3142019808292389
	pesos_i(6315) := b"1111111111111111_1111111111111111_1011100010111010_0011001000000000"; -- -0.27840888500213623
	pesos_i(6316) := b"1111111111111111_1111111111111111_1101010101111000_0001101110000000"; -- -0.16613605618476868
	pesos_i(6317) := b"0000000000000000_0000000000000000_0011001010100111_0000110011000000"; -- 0.1978614777326584
	pesos_i(6318) := b"0000000000000000_0000000000000000_0001111111001110_1000001010000000"; -- 0.12424483895301819
	pesos_i(6319) := b"0000000000000000_0000000000000000_0001001001001111_0100111111100000"; -- 0.07152270525693893
	pesos_i(6320) := b"0000000000000000_0000000000000000_0011001100100101_0101100010000000"; -- 0.19978860020637512
	pesos_i(6321) := b"1111111111111111_1111111111111111_1101000001100010_0100111011000000"; -- -0.18599994480609894
	pesos_i(6322) := b"1111111111111111_1111111111111111_1101000011000110_1010101000000000"; -- -0.18446862697601318
	pesos_i(6323) := b"0000000000000000_0000000000000000_0101001111010100_0101010000000000"; -- 0.32745862007141113
	pesos_i(6324) := b"1111111111111111_1111111111111111_1111011010000011_0010110000110000"; -- -0.03706096485257149
	pesos_i(6325) := b"0000000000000000_0000000000000000_0010100011011010_0000110100000000"; -- 0.15957719087600708
	pesos_i(6326) := b"1111111111111111_1111111111111111_1110111101010101_0111010010000000"; -- -0.06510230898857117
	pesos_i(6327) := b"0000000000000000_0000000000000000_0000000011001101_1010111001010101"; -- 0.0031384427566081285
	pesos_i(6328) := b"1111111111111111_1111111111111111_1001100011001011_1101011000000000"; -- -0.40313971042633057
	pesos_i(6329) := b"0000000000000000_0000000000000000_0011111111000110_1001001011000000"; -- 0.2491237372159958
	pesos_i(6330) := b"0000000000000000_0000000000000000_0001101111010111_1011111110000000"; -- 0.10876080393791199
	pesos_i(6331) := b"1111111111111111_1111111111111111_1111000001001110_0001111100110000"; -- -0.06130795553326607
	pesos_i(6332) := b"1111111111111111_1111111111111111_1111111110010011_0011110011100100"; -- -0.0016595786437392235
	pesos_i(6333) := b"0000000000000000_0000000000000000_0000110000010111_1101001111000000"; -- 0.04723857343196869
	pesos_i(6334) := b"0000000000000000_0000000000000000_0001011011111000_0000010011100000"; -- 0.08972197026014328
	pesos_i(6335) := b"0000000000000000_0000000000000000_0000111011010000_0011101000000000"; -- 0.05786478519439697
	pesos_i(6336) := b"1111111111111111_1111111111111111_1100100000011000_1001011011000000"; -- -0.2183748036623001
	pesos_i(6337) := b"0000000000000000_0000000000000000_0001001010011111_0011010101000000"; -- 0.07274182140827179
	pesos_i(6338) := b"0000000000000000_0000000000000000_0000010101000100_0100011101101000"; -- 0.020573103800415993
	pesos_i(6339) := b"0000000000000000_0000000000000000_0000101000001000_1100001111100000"; -- 0.03919624537229538
	pesos_i(6340) := b"0000000000000000_0000000000000000_0000100011100111_0111000010100000"; -- 0.03478149324655533
	pesos_i(6341) := b"0000000000000000_0000000000000000_0100100010100011_0110100010000000"; -- 0.28374341130256653
	pesos_i(6342) := b"1111111111111111_1111111111111111_1111101101100111_1010000100000000"; -- -0.017949998378753662
	pesos_i(6343) := b"1111111111111111_1111111111111111_1110110110001100_0011111000000000"; -- -0.07207882404327393
	pesos_i(6344) := b"1111111111111111_1111111111111111_1111010001100010_0100001101010000"; -- -0.045375626534223557
	pesos_i(6345) := b"0000000000000000_0000000000000000_0011110110010110_1111101000000000"; -- 0.24058496952056885
	pesos_i(6346) := b"1111111111111111_1111111111111111_1111000010010010_1101101111110000"; -- -0.06025910750031471
	pesos_i(6347) := b"1111111111111111_1111111111111111_1110001011110001_1011111110000000"; -- -0.11349871754646301
	pesos_i(6348) := b"0000000000000000_0000000000000000_0000110001000000_0101001000010000"; -- 0.04785645380616188
	pesos_i(6349) := b"1111111111111111_1111111111111111_1110101111001101_0011101011100000"; -- -0.07889968901872635
	pesos_i(6350) := b"0000000000000000_0000000000000000_0000110111001100_0111100000000000"; -- 0.05390119552612305
	pesos_i(6351) := b"1111111111111111_1111111111111111_1101110001011101_1011110000000000"; -- -0.13919472694396973
	pesos_i(6352) := b"1111111111111111_1111111111111111_1110010100001011_1100111101000000"; -- -0.1052885502576828
	pesos_i(6353) := b"0000000000000000_0000000000000000_0010000100111100_1011100000000000"; -- 0.12983274459838867
	pesos_i(6354) := b"1111111111111111_1111111111111111_1111010011010100_1010010011110000"; -- -0.04363030567765236
	pesos_i(6355) := b"1111111111111111_1111111111111111_1101011001111100_0010011100000000"; -- -0.16216808557510376
	pesos_i(6356) := b"0000000000000000_0000000000000000_0000111011000011_0000011011000000"; -- 0.057663366198539734
	pesos_i(6357) := b"0000000000000000_0000000000000000_0001001001111001_1101000111100000"; -- 0.07217132300138474
	pesos_i(6358) := b"0000000000000000_0000000000000000_0000001011100111_0010100010110000"; -- 0.011339705437421799
	pesos_i(6359) := b"1111111111111111_1111111111111111_1111110010100011_1001011001010100"; -- -0.013128857128322124
	pesos_i(6360) := b"0000000000000000_0000000000000000_0011000000011101_0110101100000000"; -- 0.18794888257980347
	pesos_i(6361) := b"1111111111111111_1111111111111111_1110111100011111_0101111011000000"; -- -0.06592757999897003
	pesos_i(6362) := b"0000000000000000_0000000000000000_0010000010011100_1000000110000000"; -- 0.1273880898952484
	pesos_i(6363) := b"0000000000000000_0000000000000000_0001010100110111_1010111110000000"; -- 0.08288094401359558
	pesos_i(6364) := b"1111111111111111_1111111111111111_1100111001010111_1010000111000000"; -- -0.19397534430027008
	pesos_i(6365) := b"1111111111111111_1111111111111111_1101011111100000_0110111010000000"; -- -0.15673169493675232
	pesos_i(6366) := b"1111111111111111_1111111111111111_1110110000110111_1110000011100000"; -- -0.07727236300706863
	pesos_i(6367) := b"0000000000000000_0000000000000000_0001011111010000_1010111001000000"; -- 0.09302796423435211
	pesos_i(6368) := b"0000000000000000_0000000000000000_0011001100000111_1011111110000000"; -- 0.199336975812912
	pesos_i(6369) := b"0000000000000000_0000000000000000_0001001110010101_1010111111100000"; -- 0.07650279253721237
	pesos_i(6370) := b"0000000000000000_0000000000000000_0011110110001101_0100110100000000"; -- 0.2404373288154602
	pesos_i(6371) := b"0000000000000000_0000000000000000_0011000110111000_0011000000000000"; -- 0.19421672821044922
	pesos_i(6372) := b"0000000000000000_0000000000000000_0011101000111100_1100010011000000"; -- 0.22748975455760956
	pesos_i(6373) := b"0000000000000000_0000000000000000_0010001100001000_1111001110000000"; -- 0.1368553340435028
	pesos_i(6374) := b"1111111111111111_1111111111111111_1111101001100001_1000011110000000"; -- -0.021949321031570435
	pesos_i(6375) := b"0000000000000000_0000000000000000_0101000111100000_1000100010000000"; -- 0.31983235478401184
	pesos_i(6376) := b"1111111111111111_1111111111111111_1001000001000111_0101111010000000"; -- -0.4364109933376312
	pesos_i(6377) := b"0000000000000000_0000000000000000_0000001110111010_1111100011101000"; -- 0.014571720734238625
	pesos_i(6378) := b"0000000000000000_0000000000000000_0100010001000010_1010001000000000"; -- 0.2666417360305786
	pesos_i(6379) := b"0000000000000000_0000000000000000_0000010011111000_0000001011110000"; -- 0.019409354776144028
	pesos_i(6380) := b"1111111111111111_1111111111111111_0110110101110001_0011011100000000"; -- -0.5724912285804749
	pesos_i(6381) := b"1111111111111111_1111111111111111_1110110001101110_1111001010100000"; -- -0.07643207162618637
	pesos_i(6382) := b"0000000000000000_0000000000000000_0011100011011010_0001000100000000"; -- 0.22207742929458618
	pesos_i(6383) := b"1111111111111111_1111111111111111_1101111001011101_1101001010000000"; -- -0.13138088583946228
	pesos_i(6384) := b"1111111111111111_1111111111111111_1110101000010000_0001001010000000"; -- -0.08569225668907166
	pesos_i(6385) := b"1111111111111111_1111111111111111_1101000100110111_0010100111000000"; -- -0.18275202810764313
	pesos_i(6386) := b"1111111111111111_1111111111111111_1100000001101000_0010010110000000"; -- -0.24841085076332092
	pesos_i(6387) := b"0000000000000000_0000000000000000_0001101010011000_0111111000000000"; -- 0.1038893461227417
	pesos_i(6388) := b"1111111111111111_1111111111111111_1111100100100011_1010110110111000"; -- -0.026799337938427925
	pesos_i(6389) := b"1111111111111111_1111111111111111_1101110001011100_0101011101000000"; -- -0.13921599090099335
	pesos_i(6390) := b"1111111111111111_1111111111111111_1111000010101001_0110010100110000"; -- -0.05991523340344429
	pesos_i(6391) := b"0000000000000000_0000000000000000_0011000010010011_1110100001000000"; -- 0.18975688517093658
	pesos_i(6392) := b"0000000000000000_0000000000000000_0000010111001000_1101011110110000"; -- 0.022595863789319992
	pesos_i(6393) := b"0000000000000000_0000000000000000_0000110100111101_0010100100100000"; -- 0.05171448737382889
	pesos_i(6394) := b"1111111111111111_1111111111111111_1100111100111000_1101001100000000"; -- -0.1905391812324524
	pesos_i(6395) := b"0000000000000000_0000000000000000_0000101110100110_0001110110000000"; -- 0.045503467321395874
	pesos_i(6396) := b"1111111111111111_1111111111111111_1101111100110001_0101100100000000"; -- -0.1281532645225525
	pesos_i(6397) := b"1111111111111111_1111111111111111_1101110110100000_1010110001000000"; -- -0.13426707684993744
	pesos_i(6398) := b"1111111111111111_1111111111111111_1110110100101111_0111100110000000"; -- -0.07349434494972229
	pesos_i(6399) := b"0000000000000000_0000000000000000_0011101011011101_1011110000000000"; -- 0.22994589805603027
	pesos_i(6400) := b"0000000000000000_0000000000000000_0001111101000110_0010011010100000"; -- 0.12216416746377945
	pesos_i(6401) := b"1111111111111111_1111111111111111_1111111101011101_1000001110110111"; -- -0.002479331800714135
	pesos_i(6402) := b"0000000000000000_0000000000000000_0001100000110110_1000010101100000"; -- 0.09458192437887192
	pesos_i(6403) := b"0000000000000000_0000000000000000_0001000110101000_1001111000000000"; -- 0.06897914409637451
	pesos_i(6404) := b"1111111111111111_1111111111111111_1110100100011111_1010010101100000"; -- -0.08936087042093277
	pesos_i(6405) := b"1111111111111111_1111111111111111_1100001111010101_0011001000000000"; -- -0.23502814769744873
	pesos_i(6406) := b"0000000000000000_0000000000000000_0011101111110110_0001100001000000"; -- 0.2342238575220108
	pesos_i(6407) := b"1111111111111111_1111111111111111_1101010111001110_1111111011000000"; -- -0.16481025516986847
	pesos_i(6408) := b"1111111111111111_1111111111111111_1111001011000010_0011011110110000"; -- -0.05172397568821907
	pesos_i(6409) := b"1111111111111111_1111111111111111_1111111101001100_1010111100001110"; -- -0.0027361479587852955
	pesos_i(6410) := b"1111111111111111_1111111111111111_1110001110011011_1100101001000000"; -- -0.11090408265590668
	pesos_i(6411) := b"0000000000000000_0000000000000000_0001000011101110_1010111010000000"; -- 0.0661419928073883
	pesos_i(6412) := b"1111111111111111_1111111111111111_1010101110010101_1101110010000000"; -- -0.3297445476055145
	pesos_i(6413) := b"1111111111111111_1111111111111111_1011001001010011_1100000100000000"; -- -0.30340951681137085
	pesos_i(6414) := b"0000000000000000_0000000000000000_0001110000110001_1001111001000000"; -- 0.1101321130990982
	pesos_i(6415) := b"0000000000000000_0000000000000000_0000010101111011_1011011000111000"; -- 0.021418942138552666
	pesos_i(6416) := b"1111111111111111_1111111111111111_1010110000010100_1111000110000000"; -- -0.32780542969703674
	pesos_i(6417) := b"1111111111111111_1111111111111111_1111100110110110_1110100110101000"; -- -0.0245527233928442
	pesos_i(6418) := b"0000000000000000_0000000000000000_0011110010100111_0001010010000000"; -- 0.2369244396686554
	pesos_i(6419) := b"0000000000000000_0000000000000000_0001000110001001_1000011001000000"; -- 0.0685047060251236
	pesos_i(6420) := b"0000000000000000_0000000000000000_0001001010001011_0101111100100000"; -- 0.07243914157152176
	pesos_i(6421) := b"1111111111111111_1111111111111111_1110111110000101_0011110011000000"; -- -0.0643732100725174
	pesos_i(6422) := b"0000000000000000_0000000000000000_0011110000111101_1110100010000000"; -- 0.23531964421272278
	pesos_i(6423) := b"1111111111111111_1111111111111111_1101010001011011_1110010100000000"; -- -0.17047280073165894
	pesos_i(6424) := b"1111111111111111_1111111111111111_1100100101110010_1110110011000000"; -- -0.21309013664722443
	pesos_i(6425) := b"1111111111111111_1111111111111111_1101010111100111_1001001110000000"; -- -0.16443517804145813
	pesos_i(6426) := b"0000000000000000_0000000000000000_0101000000011000_1000011100000000"; -- 0.3128742575645447
	pesos_i(6427) := b"1111111111111111_1111111111111111_1111010111011011_0110011010000000"; -- -0.03962096571922302
	pesos_i(6428) := b"0000000000000000_0000000000000000_0000011100111101_1000010011010000"; -- 0.02828245237469673
	pesos_i(6429) := b"0000000000000000_0000000000000000_0000101011110011_0100001010000000"; -- 0.042774349451065063
	pesos_i(6430) := b"0000000000000000_0000000000000000_0010101001110000_0011011111000000"; -- 0.16577480733394623
	pesos_i(6431) := b"0000000000000000_0000000000000000_0000000010101001_0000011101100110"; -- 0.0025791763328015804
	pesos_i(6432) := b"0000000000000000_0000000000000000_0000101100001000_0001101001110000"; -- 0.04309239611029625
	pesos_i(6433) := b"0000000000000000_0000000000000000_0010111010110001_1001000100000000"; -- 0.18239694833755493
	pesos_i(6434) := b"1111111111111111_1111111111111111_1111110101001000_1111000111101100"; -- -0.010605697520077229
	pesos_i(6435) := b"0000000000000000_0000000000000000_0010010000001010_0001011001000000"; -- 0.14077891409397125
	pesos_i(6436) := b"0000000000000000_0000000000000000_0001100100010011_1101010101100000"; -- 0.09795888513326645
	pesos_i(6437) := b"0000000000000000_0000000000000000_0010111100001001_0100011111000000"; -- 0.18373535573482513
	pesos_i(6438) := b"0000000000000000_0000000000000000_0001000010100010_1001111010100000"; -- 0.0649813786149025
	pesos_i(6439) := b"1111111111111111_1111111111111111_1011010000000100_0110110000000000"; -- -0.29680752754211426
	pesos_i(6440) := b"0000000000000000_0000000000000000_0111011000101001_0111101110000000"; -- 0.46157047152519226
	pesos_i(6441) := b"0000000000000000_0000000000000000_0000010110000100_1110010100111000"; -- 0.02155907265841961
	pesos_i(6442) := b"1111111111111111_1111111111111111_1100101100000111_0101110000000000"; -- -0.20691895484924316
	pesos_i(6443) := b"1111111111111111_1111111111111111_1100101100100001_0011111101000000"; -- -0.20652393996715546
	pesos_i(6444) := b"1111111111111111_1111111111111111_1100110110000000_0010100111000000"; -- -0.19726313650608063
	pesos_i(6445) := b"0000000000000000_0000000000000000_0010110011010100_1101000111000000"; -- 0.17512236535549164
	pesos_i(6446) := b"1111111111111111_1111111111111111_1100011100110010_1000100001000000"; -- -0.22188518941402435
	pesos_i(6447) := b"0000000000000000_0000000000000000_0000100111010110_1111110010110000"; -- 0.03843669220805168
	pesos_i(6448) := b"0000000000000000_0000000000000000_0011100101011100_1100001000000000"; -- 0.22407162189483643
	pesos_i(6449) := b"1111111111111111_1111111111111111_1110111111110011_1000100010100000"; -- -0.06269022077322006
	pesos_i(6450) := b"1111111111111111_1111111111111111_1101110010010100_0110111010000000"; -- -0.13836011290550232
	pesos_i(6451) := b"0000000000000000_0000000000000000_0001110011010101_1000100001000000"; -- 0.11263324320316315
	pesos_i(6452) := b"0000000000000000_0000000000000000_0010011110000101_1001100000000000"; -- 0.15438222885131836
	pesos_i(6453) := b"0000000000000000_0000000000000000_0010100000011110_0000111110000000"; -- 0.15670868754386902
	pesos_i(6454) := b"0000000000000000_0000000000000000_0001110001011001_1100100101000000"; -- 0.11074502766132355
	pesos_i(6455) := b"0000000000000000_0000000000000000_0010010101100001_0001110000000000"; -- 0.1460130214691162
	pesos_i(6456) := b"1111111111111111_1111111111111111_1100000011011111_1101100101000000"; -- -0.24658434092998505
	pesos_i(6457) := b"0000000000000000_0000000000000000_0100100111001101_1011101010000000"; -- 0.2882954180240631
	pesos_i(6458) := b"1111111111111111_1111111111111111_1100100101101000_1011101001000000"; -- -0.21324573457241058
	pesos_i(6459) := b"0000000000000000_0000000000000000_0011001011000111_1010001010000000"; -- 0.1983586847782135
	pesos_i(6460) := b"0000000000000000_0000000000000000_0010101111111001_1111111100000000"; -- 0.17178338766098022
	pesos_i(6461) := b"1111111111111111_1111111111111111_1101010000110110_0001010001000000"; -- -0.1710498183965683
	pesos_i(6462) := b"1111111111111111_1111111111111111_1110001111010000_0101100101100000"; -- -0.1101020947098732
	pesos_i(6463) := b"0000000000000000_0000000000000000_0011001111000101_1101010010000000"; -- 0.20223739743232727
	pesos_i(6464) := b"0000000000000000_0000000000000000_0011000010111010_0001010000000000"; -- 0.1903393268585205
	pesos_i(6465) := b"0000000000000000_0000000000000000_0001100010110100_1001011000100000"; -- 0.0965055301785469
	pesos_i(6466) := b"0000000000000000_0000000000000000_0001001100011101_1111000110100000"; -- 0.07467565685510635
	pesos_i(6467) := b"0000000000000000_0000000000000000_0100011001001110_0100111110000000"; -- 0.27463242411613464
	pesos_i(6468) := b"0000000000000000_0000000000000000_0001101011010000_1011111011100000"; -- 0.1047477051615715
	pesos_i(6469) := b"0000000000000000_0000000000000000_0001000110001001_0100000000000000"; -- 0.06850051879882812
	pesos_i(6470) := b"0000000000000000_0000000000000000_0101111111100111_0010100010000000"; -- 0.3746209442615509
	pesos_i(6471) := b"0000000000000000_0000000000000000_0000011011010000_0110101100001000"; -- 0.026617707684636116
	pesos_i(6472) := b"0000000000000000_0000000000000000_0100000100011000_0111000010000000"; -- 0.25427916646003723
	pesos_i(6473) := b"0000000000000000_0000000000000000_0001001010010100_1110100011000000"; -- 0.07258467376232147
	pesos_i(6474) := b"0000000000000000_0000000000000000_0010011101110101_0001110110000000"; -- 0.15413078665733337
	pesos_i(6475) := b"1111111111111111_1111111111111111_1110000101100101_1011011111100000"; -- -0.11954165250062943
	pesos_i(6476) := b"0000000000000000_0000000000000000_0010001110010110_1010010001000000"; -- 0.13901735842227936
	pesos_i(6477) := b"0000000000000000_0000000000000000_0001111011101100_0011111110100000"; -- 0.12079236656427383
	pesos_i(6478) := b"1111111111111111_1111111111111111_1011101011001001_1111111010000000"; -- -0.27035531401634216
	pesos_i(6479) := b"0000000000000000_0000000000000000_0001010001000111_0000001010100000"; -- 0.07920853048563004
	pesos_i(6480) := b"0000000000000000_0000000000000000_0000110011010111_1111010100010000"; -- 0.05017024651169777
	pesos_i(6481) := b"0000000000000000_0000000000000000_0110111001110010_0111100010000000"; -- 0.43143418431282043
	pesos_i(6482) := b"1111111111111111_1111111111111111_1111011100110100_0101011111100000"; -- -0.03435755521059036
	pesos_i(6483) := b"0000000000000000_0000000000000000_0010011011111101_0010000100000000"; -- 0.1522999405860901
	pesos_i(6484) := b"0000000000000000_0000000000000000_0010110101011110_0101111010000000"; -- 0.17722120881080627
	pesos_i(6485) := b"1111111111111111_1111111111111111_1111100001110111_0000001100111000"; -- -0.02943401224911213
	pesos_i(6486) := b"0000000000000000_0000000000000000_0011011000000100_0011000000000000"; -- 0.21100139617919922
	pesos_i(6487) := b"0000000000000000_0000000000000000_0011011011101011_0111100111000000"; -- 0.2145305722951889
	pesos_i(6488) := b"0000000000000000_0000000000000000_0010010010100001_1110110001000000"; -- 0.14309574663639069
	pesos_i(6489) := b"0000000000000000_0000000000000000_0100001101000100_0010011100000000"; -- 0.26275867223739624
	pesos_i(6490) := b"1111111111111111_1111111111111111_1111001100010100_1110000100000000"; -- -0.05046266317367554
	pesos_i(6491) := b"1111111111111111_1111111111111111_1011111100001110_0101111110000000"; -- -0.25368693470954895
	pesos_i(6492) := b"0000000000000000_0000000000000000_0001000111011001_0110100110100000"; -- 0.0697237029671669
	pesos_i(6493) := b"1111111111111111_1111111111111111_1111011100110100_0001001100000000"; -- -0.03436166048049927
	pesos_i(6494) := b"1111111111111111_1111111111111111_1111000000011000_0111101110100000"; -- -0.06212642043828964
	pesos_i(6495) := b"1111111111111111_1111111111111111_1111000001011011_1011010010010000"; -- -0.061100687831640244
	pesos_i(6496) := b"1111111111111111_1111111111111111_1100000001111110_1001000110000000"; -- -0.24806872010231018
	pesos_i(6497) := b"0000000000000000_0000000000000000_0000010001010010_1100110110111000"; -- 0.016888482496142387
	pesos_i(6498) := b"0000000000000000_0000000000000000_0010011011011000_0010000000000000"; -- 0.1517353057861328
	pesos_i(6499) := b"0000000000000000_0000000000000000_0100011110011101_0111111010000000"; -- 0.2797469198703766
	pesos_i(6500) := b"0000000000000000_0000000000000000_0001100100111011_1000111010000000"; -- 0.098565012216568
	pesos_i(6501) := b"0000000000000000_0000000000000000_0011001000101000_1011011000000000"; -- 0.19593369960784912
	pesos_i(6502) := b"0000000000000000_0000000000000000_0001100111111110_1001101011100000"; -- 0.10154121369123459
	pesos_i(6503) := b"0000000000000000_0000000000000000_0101011110000110_0100010100000000"; -- 0.3418925404548645
	pesos_i(6504) := b"1111111111111111_1111111111111111_1111101000100100_1100100101111000"; -- -0.022876175120472908
	pesos_i(6505) := b"0000000000000000_0000000000000000_0000000011010010_1000000100110011"; -- 0.0032120465766638517
	pesos_i(6506) := b"0000000000000000_0000000000000000_0110100110000000_1001011110000000"; -- 0.41211840510368347
	pesos_i(6507) := b"0000000000000000_0000000000000000_0100100010100001_0101101000000000"; -- 0.2837120294570923
	pesos_i(6508) := b"1111111111111111_1111111111111111_1110000000000011_1110110101000000"; -- -0.12494008243083954
	pesos_i(6509) := b"0000000000000000_0000000000000000_0010010110111000_0101100000000000"; -- 0.14734411239624023
	pesos_i(6510) := b"0000000000000000_0000000000000000_0100001001011010_0010001110000000"; -- 0.2591879069805145
	pesos_i(6511) := b"0000000000000000_0000000000000000_0001100000111111_1010000000000000"; -- 0.09472084045410156
	pesos_i(6512) := b"1111111111111111_1111111111111111_1100000000000111_0001000111000000"; -- -0.24989213049411774
	pesos_i(6513) := b"1111111111111111_1111111111111111_1010111000000000_0111100110000000"; -- -0.3203052580356598
	pesos_i(6514) := b"0000000000000000_0000000000000000_0000001100011010_0111010100001000"; -- 0.01212245412170887
	pesos_i(6515) := b"1111111111111111_1111111111111111_1101100010011000_1010001100000000"; -- -0.1539209485054016
	pesos_i(6516) := b"0000000000000000_0000000000000000_0001100111101000_0110100011000000"; -- 0.10120253264904022
	pesos_i(6517) := b"1111111111111111_1111111111111111_1001010101110101_0100100100000000"; -- -0.4161791205406189
	pesos_i(6518) := b"1111111111111111_1111111111111111_1111111010100010_0100001000001100"; -- -0.0053366394713521
	pesos_i(6519) := b"0000000000000000_0000000000000000_0011001110010110_1100000100000000"; -- 0.20151907205581665
	pesos_i(6520) := b"1111111111111111_1111111111111111_1110000111100100_1001000001000000"; -- -0.11760614812374115
	pesos_i(6521) := b"0000000000000000_0000000000000000_0010100110110110_1101011011000000"; -- 0.16294614970684052
	pesos_i(6522) := b"1111111111111111_1111111111111111_1111111100010000_1100001110101001"; -- -0.0036504471208900213
	pesos_i(6523) := b"1111111111111111_1111111111111111_1101001100000111_0110011100000000"; -- -0.17566829919815063
	pesos_i(6524) := b"1111111111111111_1111111111111111_1111000011011000_1101101000110000"; -- -0.05919109657406807
	pesos_i(6525) := b"1111111111111111_1111111111111111_1110000101101111_0110011100100000"; -- -0.11939387768507004
	pesos_i(6526) := b"0000000000000000_0000000000000000_0000001001011110_1110110001011100"; -- 0.009260914288461208
	pesos_i(6527) := b"0000000000000000_0000000000000000_0100011100100101_0011111010000000"; -- 0.27791205048561096
	pesos_i(6528) := b"0000000000000000_0000000000000000_0000010100011111_0110011100010000"; -- 0.020010415464639664
	pesos_i(6529) := b"1111111111111111_1111111111111111_1110101011011100_0110111011100000"; -- -0.08257395774126053
	pesos_i(6530) := b"0000000000000000_0000000000000000_0100011110100111_0101110010000000"; -- 0.2798974812030792
	pesos_i(6531) := b"1111111111111111_1111111111111111_1111011001001100_1000111100110000"; -- -0.037894297391176224
	pesos_i(6532) := b"0000000000000000_0000000000000000_0001000001011111_1110100101000000"; -- 0.06396348774433136
	pesos_i(6533) := b"1111111111111111_1111111111111111_1011001110011001_1011101000000000"; -- -0.2984355688095093
	pesos_i(6534) := b"0000000000000000_0000000000000000_0110110010011000_0101001000000000"; -- 0.4241992235183716
	pesos_i(6535) := b"0000000000000000_0000000000000000_0001000111100111_1001001010000000"; -- 0.0699397623538971
	pesos_i(6536) := b"1111111111111111_1111111111111111_1110111110101010_0011100110100000"; -- -0.06380882114171982
	pesos_i(6537) := b"0000000000000000_0000000000000000_0010110001111010_0011110110000000"; -- 0.1737402379512787
	pesos_i(6538) := b"0000000000000000_0000000000000000_0010010011110111_1010001011000000"; -- 0.1444036215543747
	pesos_i(6539) := b"0000000000000000_0000000000000000_0001111010011100_0110101111100000"; -- 0.11957430094480515
	pesos_i(6540) := b"0000000000000000_0000000000000000_0010011011000001_0001101100000000"; -- 0.15138405561447144
	pesos_i(6541) := b"1111111111111111_1111111111111111_1101001111001011_1101111001000000"; -- -0.17267046868801117
	pesos_i(6542) := b"0000000000000000_0000000000000000_0101010010100001_1100011010000000"; -- 0.3305934965610504
	pesos_i(6543) := b"0000000000000000_0000000000000000_0000111100111100_0011111001110000"; -- 0.05951299890875816
	pesos_i(6544) := b"1111111111111111_1111111111111111_1011110101011010_1110101100000000"; -- -0.2603314518928528
	pesos_i(6545) := b"0000000000000000_0000000000000000_0111101101000001_0001100110000000"; -- 0.4814620912075043
	pesos_i(6546) := b"0000000000000000_0000000000000000_0011101011001001_1101010010000000"; -- 0.22964218258857727
	pesos_i(6547) := b"0000000000000000_0000000000000000_0100010110101101_0010001110000000"; -- 0.272173136472702
	pesos_i(6548) := b"0000000000000000_0000000000000000_0011110000001010_1101001100000000"; -- 0.2345401644706726
	pesos_i(6549) := b"1111111111111111_1111111111111111_1101001011100111_0110111110000000"; -- -0.17615607380867004
	pesos_i(6550) := b"0000000000000000_0000000000000000_0011100000111000_0100111000000000"; -- 0.21960914134979248
	pesos_i(6551) := b"1111111111111111_1111111111111111_1011011110110100_1111001100000000"; -- -0.2823951840400696
	pesos_i(6552) := b"1111111111111111_1111111111111111_1010001011101100_1000100110000000"; -- -0.3635782301425934
	pesos_i(6553) := b"1111111111111111_1111111111111111_1111110001101110_1000001000001100"; -- -0.013938781805336475
	pesos_i(6554) := b"0000000000000000_0000000000000000_0010000010110011_1011110100000000"; -- 0.12774258852005005
	pesos_i(6555) := b"0000000000000000_0000000000000000_0110110100000000_1010010000000000"; -- 0.42579102516174316
	pesos_i(6556) := b"1111111111111111_1111111111111111_1111100101101001_1101100101000000"; -- -0.025728628039360046
	pesos_i(6557) := b"0000000000000000_0000000000000000_0011100000010110_0101101100000000"; -- 0.21909111738204956
	pesos_i(6558) := b"0000000000000000_0000000000000000_0000100000100111_0000010001000000"; -- 0.031845346093177795
	pesos_i(6559) := b"0000000000000000_0000000000000000_0010010100101010_1001000010000000"; -- 0.14518073201179504
	pesos_i(6560) := b"1111111111111111_1111111111111111_1101011001000110_0100011001000000"; -- -0.16299019753932953
	pesos_i(6561) := b"1111111111111111_1111111111111111_1111011111101100_1111010101000000"; -- -0.031540557742118835
	pesos_i(6562) := b"0000000000000000_0000000000000000_0100111100000100_1111100100000000"; -- 0.3086696267127991
	pesos_i(6563) := b"0000000000000000_0000000000000000_0010011010110100_0100011011000000"; -- 0.15118829905986786
	pesos_i(6564) := b"0000000000000000_0000000000000000_0101010101010010_0101010010000000"; -- 0.3332875072956085
	pesos_i(6565) := b"0000000000000000_0000000000000000_0011001011011111_1101100101000000"; -- 0.19872815907001495
	pesos_i(6566) := b"0000000000000000_0000000000000000_0010010111010111_0000010010000000"; -- 0.147812157869339
	pesos_i(6567) := b"1111111111111111_1111111111111111_1111010011011101_0000110101100000"; -- -0.04350201040506363
	pesos_i(6568) := b"0000000000000000_0000000000000000_1001010001010011_1101011000000000"; -- 0.5794042348861694
	pesos_i(6569) := b"0000000000000000_0000000000000000_0101111100010110_0110010100000000"; -- 0.3714354634284973
	pesos_i(6570) := b"0000000000000000_0000000000000000_0101101010101001_1110000100000000"; -- 0.35415464639663696
	pesos_i(6571) := b"0000000000000000_0000000000000000_0000000000110110_1010110001010011"; -- 0.0008342458750121295
	pesos_i(6572) := b"0000000000000000_0000000000000000_0000001100010101_1011100011110000"; -- 0.012050207704305649
	pesos_i(6573) := b"0000000000000000_0000000000000000_0110010000100111_1011011110000000"; -- 0.3912310302257538
	pesos_i(6574) := b"1111111111111111_1111111111111111_1001111010110010_1111010100000000"; -- -0.38008183240890503
	pesos_i(6575) := b"0000000000000000_0000000000000000_0011111011001010_1010001001000000"; -- 0.2452794462442398
	pesos_i(6576) := b"0000000000000000_0000000000000000_1000011110000010_1011010100000000"; -- 0.5293381810188293
	pesos_i(6577) := b"1111111111111111_1111111111111111_1111010100100101_0110110110110000"; -- -0.0423976369202137
	pesos_i(6578) := b"0000000000000000_0000000000000000_0010010011101101_1011010010000000"; -- 0.14425209164619446
	pesos_i(6579) := b"0000000000000000_0000000000000000_0000101101101100_0001001011000000"; -- 0.04461781680583954
	pesos_i(6580) := b"0000000000000000_0000000000000000_0010001010101010_1101100010000000"; -- 0.13541939854621887
	pesos_i(6581) := b"0000000000000000_0000000000000000_0100000000010111_1110011100000000"; -- 0.2503647208213806
	pesos_i(6582) := b"0000000000000000_0000000000000000_0101001010011110_1011000000000000"; -- 0.32273387908935547
	pesos_i(6583) := b"1111111111111111_1111111111111111_1111001000010011_1010110110100000"; -- -0.05438723415136337
	pesos_i(6584) := b"1111111111111111_1111111111111111_1111110000110010_1111000011101000"; -- -0.014847701415419579
	pesos_i(6585) := b"1111111111111111_1111111111111111_1111101101111010_1111000000001000"; -- -0.017655370756983757
	pesos_i(6586) := b"0000000000000000_0000000000000000_0001001110010111_1000100111000000"; -- 0.07653103768825531
	pesos_i(6587) := b"0000000000000000_0000000000000000_0110011001001010_1000011100000000"; -- 0.3995746970176697
	pesos_i(6588) := b"0000000000000000_0000000000000000_0001000001100000_1011111011000000"; -- 0.0639762133359909
	pesos_i(6589) := b"1111111111111111_1111111111111111_1100111100100011_1110010010000000"; -- -0.19085857272148132
	pesos_i(6590) := b"0000000000000000_0000000000000000_0010010101111000_1110110100000000"; -- 0.14637643098831177
	pesos_i(6591) := b"0000000000000000_0000000000000000_0011001001010101_1010000110000000"; -- 0.19661912322044373
	pesos_i(6592) := b"1111111111111111_1111111111111111_1100111111011100_0110100111000000"; -- -0.188043013215065
	pesos_i(6593) := b"0000000000000000_0000000000000000_0000001000001010_0001011001000000"; -- 0.007966414093971252
	pesos_i(6594) := b"1111111111111111_1111111111111111_1111111001011001_0111010010111100"; -- -0.006447509862482548
	pesos_i(6595) := b"0000000000000000_0000000000000000_0011101111110010_1010010001000000"; -- 0.23417116701602936
	pesos_i(6596) := b"1111111111111111_1111111111111111_1100111100011101_1101111010000000"; -- -0.19095048308372498
	pesos_i(6597) := b"0000000000000000_0000000000000000_0000011001110110_1101100110111000"; -- 0.025251014158129692
	pesos_i(6598) := b"0000000000000000_0000000000000000_0100001101100001_0011000000000000"; -- 0.2632017135620117
	pesos_i(6599) := b"1111111111111111_1111111111111111_1110111001011101_1000110000100000"; -- -0.06888508051633835
	pesos_i(6600) := b"0000000000000000_0000000000000000_0010010000100111_0100000010000000"; -- 0.1412239372730255
	pesos_i(6601) := b"0000000000000000_0000000000000000_0100111110000100_0001000010000000"; -- 0.3106088936328888
	pesos_i(6602) := b"1111111111111111_1111111111111111_1110100111110000_0010101001000000"; -- -0.08617912232875824
	pesos_i(6603) := b"0000000000000000_0000000000000000_0011010101001000_1110110101000000"; -- 0.20814402401447296
	pesos_i(6604) := b"0000000000000000_0000000000000000_0101011011111001_0001111100000000"; -- 0.33973878622055054
	pesos_i(6605) := b"0000000000000000_0000000000000000_0010000101000011_1011010111000000"; -- 0.12993942201137543
	pesos_i(6606) := b"1111111111111111_1111111111111111_1111100000010101_0001111101111000"; -- -0.030927689746022224
	pesos_i(6607) := b"0000000000000000_0000000000000000_0100110100110111_0001111000000000"; -- 0.30162227153778076
	pesos_i(6608) := b"1111111111111111_1111111111111111_1010011010011000_1100110100000000"; -- -0.34923094511032104
	pesos_i(6609) := b"0000000000000000_0000000000000000_0000101111010011_1111000111000000"; -- 0.04620276391506195
	pesos_i(6610) := b"0000000000000000_0000000000000000_0000101000111000_1110101011000000"; -- 0.03993098437786102
	pesos_i(6611) := b"0000000000000000_0000000000000000_0001111000110000_0110110100000000"; -- 0.11792641878128052
	pesos_i(6612) := b"0000000000000000_0000000000000000_0001001011101110_1101100011100000"; -- 0.07395701855421066
	pesos_i(6613) := b"1111111111111111_1111111111111111_1101110100000100_0100001100000000"; -- -0.13665372133255005
	pesos_i(6614) := b"1111111111111111_1111111111111111_1100111111100000_0010011010000000"; -- -0.18798598647117615
	pesos_i(6615) := b"0000000000000000_0000000000000000_0110010011110101_0101000110000000"; -- 0.3943682610988617
	pesos_i(6616) := b"0000000000000000_0000000000000000_0000100100111100_0001111011100000"; -- 0.03607361763715744
	pesos_i(6617) := b"0000000000000000_0000000000000000_0101100100110001_1011101100000000"; -- 0.3484150767326355
	pesos_i(6618) := b"1111111111111111_1111111111111111_1100101111100001_1001110000000000"; -- -0.20358872413635254
	pesos_i(6619) := b"1111111111111111_1111111111111111_1110100101101011_0101111010000000"; -- -0.08820542693138123
	pesos_i(6620) := b"0000000000000000_0000000000000000_0001001110000011_1011001000000000"; -- 0.07622826099395752
	pesos_i(6621) := b"1111111111111111_1111111111111111_1110000101001100_1000101111100000"; -- -0.11992574483156204
	pesos_i(6622) := b"0000000000000000_0000000000000000_0001000000111100_1011001000100000"; -- 0.06342614442110062
	pesos_i(6623) := b"0000000000000000_0000000000000000_0000110010101100_1001011111010000"; -- 0.049508560448884964
	pesos_i(6624) := b"1111111111111111_1111111111111111_1101000001011100_1011010010000000"; -- -0.18608543276786804
	pesos_i(6625) := b"1111111111111111_1111111111111111_1111101000001011_1101100011100000"; -- -0.023256726562976837
	pesos_i(6626) := b"1111111111111111_1111111111111111_1110111110000010_0100001111100000"; -- -0.06441856175661087
	pesos_i(6627) := b"0000000000000000_0000000000000000_0100100011001001_0011111000000000"; -- 0.2843207120895386
	pesos_i(6628) := b"0000000000000000_0000000000000000_0010111111101011_1100110010000000"; -- 0.18719175457954407
	pesos_i(6629) := b"0000000000000000_0000000000000000_0101110001110000_1010010010000000"; -- 0.36109378933906555
	pesos_i(6630) := b"0000000000000000_0000000000000000_0001010100111111_0011111000100000"; -- 0.08299625664949417
	pesos_i(6631) := b"0000000000000000_0000000000000000_0010000101010101_1111010100000000"; -- 0.13021785020828247
	pesos_i(6632) := b"1111111111111111_1111111111111111_1100001111111100_0100011011000000"; -- -0.23443181812763214
	pesos_i(6633) := b"0000000000000000_0000000000000000_0100000001010100_1110110010000000"; -- 0.2512958347797394
	pesos_i(6634) := b"0000000000000000_0000000000000000_0110000110011111_1011111010000000"; -- 0.3813437521457672
	pesos_i(6635) := b"0000000000000000_0000000000000000_0101110100001011_0011011000000000"; -- 0.36345231533050537
	pesos_i(6636) := b"0000000000000000_0000000000000000_0001100101111101_1000100010100000"; -- 0.09957174211740494
	pesos_i(6637) := b"0000000000000000_0000000000000000_0000101011010000_0000011100100000"; -- 0.042236752808094025
	pesos_i(6638) := b"0000000000000000_0000000000000000_0111011001110111_1101001100000000"; -- 0.4627658724784851
	pesos_i(6639) := b"0000000000000000_0000000000000000_0011110110101010_1010000100000000"; -- 0.24088484048843384
	pesos_i(6640) := b"0000000000000000_0000000000000000_0000011001111101_1110101000111000"; -- 0.025358809158205986
	pesos_i(6641) := b"1111111111111111_1111111111111111_1010110101000111_1011010100000000"; -- -0.32312458753585815
	pesos_i(6642) := b"1111111111111111_1111111111111111_1111111000011001_0010101001001000"; -- -0.0074285101145505905
	pesos_i(6643) := b"1111111111111111_1111111111111111_1010001101100001_1011111000000000"; -- -0.3617898225784302
	pesos_i(6644) := b"1111111111111111_1111111111111111_1110000100000011_0110111101000000"; -- -0.12104134261608124
	pesos_i(6645) := b"1111111111111111_1111111111111111_1001000101011110_0001101000000000"; -- -0.43215787410736084
	pesos_i(6646) := b"1111111111111111_1111111111111111_1001000110100001_0010111110000000"; -- -0.43113425374031067
	pesos_i(6647) := b"0000000000000000_0000000000000000_0001100010100010_1000010100100000"; -- 0.09622985869646072
	pesos_i(6648) := b"1111111111111111_1111111111111111_1110101100100111_0111100011000000"; -- -0.08142895996570587
	pesos_i(6649) := b"0000000000000000_0000000000000000_0011100111111111_1100101110000000"; -- 0.2265593707561493
	pesos_i(6650) := b"1111111111111111_1111111111111111_1110111001000100_1110100000000000"; -- -0.06926107406616211
	pesos_i(6651) := b"1111111111111111_1111111111111111_1100110000000100_1110101110000000"; -- -0.2030499279499054
	pesos_i(6652) := b"0000000000000000_0000000000000000_0110000101111111_1100000000000000"; -- 0.3808555603027344
	pesos_i(6653) := b"0000000000000000_0000000000000000_0001110100110110_0101100010100000"; -- 0.11411050707101822
	pesos_i(6654) := b"0000000000000000_0000000000000000_0000001111101001_0101001110000000"; -- 0.015279024839401245
	pesos_i(6655) := b"0000000000000000_0000000000000000_0000101011000111_0010010110000000"; -- 0.04210123419761658
	pesos_i(6656) := b"0000000000000000_0000000000000000_0000011010001100_0101010101001000"; -- 0.02557881362736225
	pesos_i(6657) := b"0000000000000000_0000000000000000_0000010101000110_1000101010011000"; -- 0.02060762606561184
	pesos_i(6658) := b"0000000000000000_0000000000000000_0011011011000100_0000001011000000"; -- 0.21392838656902313
	pesos_i(6659) := b"0000000000000000_0000000000000000_0001101011001010_0100110110000000"; -- 0.10464939475059509
	pesos_i(6660) := b"0000000000000000_0000000000000000_0000010001100011_1010011111000000"; -- 0.017145618796348572
	pesos_i(6661) := b"1111111111111111_1111111111111111_1001000000001000_0101110010000000"; -- -0.4373724162578583
	pesos_i(6662) := b"0000000000000000_0000000000000000_0001101000011100_1001110010100000"; -- 0.10199908167123795
	pesos_i(6663) := b"0000000000000000_0000000000000000_0000011001101001_0010111010100000"; -- 0.025042451918125153
	pesos_i(6664) := b"0000000000000000_0000000000000000_0110000110011111_1111001110000000"; -- 0.3813469111919403
	pesos_i(6665) := b"0000000000000000_0000000000000000_0010111101111111_1111011100000000"; -- 0.18554633855819702
	pesos_i(6666) := b"0000000000000000_0000000000000000_0100101101100010_0011000110000000"; -- 0.2944670617580414
	pesos_i(6667) := b"0000000000000000_0000000000000000_0000000101011000_1101111011000100"; -- 0.005262301303446293
	pesos_i(6668) := b"0000000000000000_0000000000000000_0011101001010111_1000011110000000"; -- 0.22789809107780457
	pesos_i(6669) := b"1111111111111111_1111111111111111_1111011110000110_1110001100110000"; -- -0.03309803083539009
	pesos_i(6670) := b"1111111111111111_1111111111111111_1110001110011111_0010010100000000"; -- -0.11085289716720581
	pesos_i(6671) := b"0000000000000000_0000000000000000_0000100000110111_1101100110000000"; -- 0.03210219740867615
	pesos_i(6672) := b"1111111111111111_1111111111111111_1111000101000001_0100100101000000"; -- -0.0575975626707077
	pesos_i(6673) := b"0000000000000000_0000000000000000_0101001011001110_1100011100000000"; -- 0.3234676718711853
	pesos_i(6674) := b"1111111111111111_1111111111111111_1111011101011010_0000011000010000"; -- -0.03378259763121605
	pesos_i(6675) := b"1111111111111111_1111111111111111_1100110010101111_1010010010000000"; -- -0.20044490694999695
	pesos_i(6676) := b"0000000000000000_0000000000000000_0101000110010111_0111000000000000"; -- 0.31871700286865234
	pesos_i(6677) := b"1111111111111111_1111111111111111_1110010011101111_0001001000000000"; -- -0.10572707653045654
	pesos_i(6678) := b"0000000000000000_0000000000000000_0110110101110100_0111010000000000"; -- 0.42755818367004395
	pesos_i(6679) := b"0000000000000000_0000000000000000_0000110011110110_1110000001000000"; -- 0.05064202845096588
	pesos_i(6680) := b"1111111111111111_1111111111111111_1011101111101111_0000100110000000"; -- -0.26588383316993713
	pesos_i(6681) := b"1111111111111111_1111111111111111_1111010011101110_0010001110010000"; -- -0.043241288512945175
	pesos_i(6682) := b"0000000000000000_0000000000000000_0001101011101110_1101000111100000"; -- 0.10520660132169724
	pesos_i(6683) := b"1111111111111111_1111111111111111_1101110000111000_1000100010000000"; -- -0.13976237177848816
	pesos_i(6684) := b"1111111111111111_1111111111111111_1111010100100000_1010011100110000"; -- -0.042470503598451614
	pesos_i(6685) := b"0000000000000000_0000000000000000_0011010000010110_0011000101000000"; -- 0.2034636288881302
	pesos_i(6686) := b"1111111111111111_1111111111111111_1111111100111110_0010100100010111"; -- -0.002957755932584405
	pesos_i(6687) := b"0000000000000000_0000000000000000_0011001100101000_1011011010000000"; -- 0.1998399794101715
	pesos_i(6688) := b"0000000000000000_0000000000000000_0000001111110001_1110100101101100"; -- 0.01541003119200468
	pesos_i(6689) := b"0000000000000000_0000000000000000_0011110010010100_0001110101000000"; -- 0.23663504421710968
	pesos_i(6690) := b"0000000000000000_0000000000000000_0010111101110011_1100111101000000"; -- 0.1853608638048172
	pesos_i(6691) := b"0000000000000000_0000000000000000_0010100011000001_0111001010000000"; -- 0.15920177102088928
	pesos_i(6692) := b"0000000000000000_0000000000000000_0001111000101001_1111010010000000"; -- 0.11782768368721008
	pesos_i(6693) := b"0000000000000000_0000000000000000_0010110110101010_0111010101000000"; -- 0.17838223278522491
	pesos_i(6694) := b"0000000000000000_0000000000000000_0001111001101100_0100010000100000"; -- 0.11883950978517532
	pesos_i(6695) := b"0000000000000000_0000000000000000_0101101010101010_0000001000000000"; -- 0.35415661334991455
	pesos_i(6696) := b"0000000000000000_0000000000000000_0101111100010110_0100101000000000"; -- 0.3714338541030884
	pesos_i(6697) := b"0000000000000000_0000000000000000_0011001001010001_0110101011000000"; -- 0.19655482470989227
	pesos_i(6698) := b"0000000000000000_0000000000000000_0101100100011001_1011110110000000"; -- 0.34804901480674744
	pesos_i(6699) := b"1111111111111111_1111111111111111_1110101011111110_0101111011100000"; -- -0.08205611258745193
	pesos_i(6700) := b"1111111111111111_1111111111111111_1101000000010000_1011110010000000"; -- -0.18724462389945984
	pesos_i(6701) := b"0000000000000000_0000000000000000_0010100010110101_1111010011000000"; -- 0.15902642905712128
	pesos_i(6702) := b"1111111111111111_1111111111111111_1110011001000111_1011011000000000"; -- -0.10046827793121338
	pesos_i(6703) := b"0000000000000000_0000000000000000_0101110001010111_1110010110000000"; -- 0.36071619391441345
	pesos_i(6704) := b"0000000000000000_0000000000000000_0100011111101011_0011010110000000"; -- 0.280932754278183
	pesos_i(6705) := b"1111111111111111_1111111111111111_1110000010010000_1101011111100000"; -- -0.12278986722230911
	pesos_i(6706) := b"1111111111111111_1111111111111111_1111100001100000_1000001110001000"; -- -0.029777316376566887
	pesos_i(6707) := b"1111111111111111_1111111111111111_1110100111111001_0111101111100000"; -- -0.08603692799806595
	pesos_i(6708) := b"1111111111111111_1111111111111111_1110111001011011_1011111001000000"; -- -0.06891261041164398
	pesos_i(6709) := b"0000000000000000_0000000000000000_0000100010110001_0001011001000000"; -- 0.03395213186740875
	pesos_i(6710) := b"0000000000000000_0000000000000000_0111111011110000_1101000010000000"; -- 0.49586203694343567
	pesos_i(6711) := b"1111111111111111_1111111111111111_1101100111110110_0011001011000000"; -- -0.14858706295490265
	pesos_i(6712) := b"0000000000000000_0000000000000000_0011100111111101_0011100011000000"; -- 0.2265201061964035
	pesos_i(6713) := b"0000000000000000_0000000000000000_0011000101101100_0101100100000000"; -- 0.193059504032135
	pesos_i(6714) := b"1111111111111111_1111111111111111_1110101100011000_0110011000100000"; -- -0.08165895193815231
	pesos_i(6715) := b"0000000000000000_0000000000000000_0011001010001010_0101101110000000"; -- 0.19742366671562195
	pesos_i(6716) := b"1111111111111111_1111111111111111_1111111100100100_1110010110011011"; -- -0.003343248041346669
	pesos_i(6717) := b"0000000000000000_0000000000000000_0010011101110101_1101010011000000"; -- 0.15414170920848846
	pesos_i(6718) := b"1111111111111111_1111111111111111_1110101100110001_1101110010000000"; -- -0.08127042651176453
	pesos_i(6719) := b"1111111111111111_1111111111111111_1111101010000011_1011111001011000"; -- -0.021427253261208534
	pesos_i(6720) := b"0000000000000000_0000000000000000_0000101111111000_0110001110100000"; -- 0.04675886780023575
	pesos_i(6721) := b"1111111111111111_1111111111111111_1010001100011000_1000001000000000"; -- -0.3629072904586792
	pesos_i(6722) := b"0000000000000000_0000000000000000_0000101010111010_0011001000000000"; -- 0.04190361499786377
	pesos_i(6723) := b"0000000000000000_0000000000000000_0010010110101011_1101110010000000"; -- 0.14715364575386047
	pesos_i(6724) := b"0000000000000000_0000000000000000_0100000100101011_0011000100000000"; -- 0.2545652985572815
	pesos_i(6725) := b"0000000000000000_0000000000000000_0000100010010000_1110000101000000"; -- 0.03346069157123566
	pesos_i(6726) := b"1111111111111111_1111111111111111_1010000011110001_0001100010000000"; -- -0.3713211715221405
	pesos_i(6727) := b"1111111111111111_1111111111111111_1011101001011011_0111011000000000"; -- -0.272041916847229
	pesos_i(6728) := b"1111111111111111_1111111111111111_1110000110110100_0000111001100000"; -- -0.11834631115198135
	pesos_i(6729) := b"0000000000000000_0000000000000000_0011011101111011_0000101011000000"; -- 0.21672122180461884
	pesos_i(6730) := b"1111111111111111_1111111111111111_1001011100010110_0101111010000000"; -- -0.4098149240016937
	pesos_i(6731) := b"0000000000000000_0000000000000000_0101100101001100_1000010110000000"; -- 0.3488238751888275
	pesos_i(6732) := b"0000000000000000_0000000000000000_0101100100110110_0001101000000000"; -- 0.34848177433013916
	pesos_i(6733) := b"1111111111111111_1111111111111111_1101000010110011_0100011011000000"; -- -0.18476445972919464
	pesos_i(6734) := b"0000000000000000_0000000000000000_0011010011110000_1001110100000000"; -- 0.20679646730422974
	pesos_i(6735) := b"1111111111111111_1111111111111111_1110101111011011_1010011010100000"; -- -0.0786796435713768
	pesos_i(6736) := b"1111111111111111_1111111111111111_0110000110011010_1011011100000000"; -- -0.6187329888343811
	pesos_i(6737) := b"1111111111111111_1111111111111111_1110111100000110_0001111001100000"; -- -0.06631288677453995
	pesos_i(6738) := b"0000000000000000_0000000000000000_0011010101110010_1010110011000000"; -- 0.20878104865550995
	pesos_i(6739) := b"0000000000000000_0000000000000000_0011000101010110_0100010110000000"; -- 0.1927226483821869
	pesos_i(6740) := b"0000000000000000_0000000000000000_0100000110111011_1011111110000000"; -- 0.256771057844162
	pesos_i(6741) := b"0000000000000000_0000000000000000_0011011001000000_1110010011000000"; -- 0.21192769706249237
	pesos_i(6742) := b"1111111111111111_1111111111111111_1110001011100110_0111101100000000"; -- -0.11367064714431763
	pesos_i(6743) := b"0000000000000000_0000000000000000_0100001011010100_1110101100000000"; -- 0.2610613703727722
	pesos_i(6744) := b"0000000000000000_0000000000000000_0001001000100111_0010100011000000"; -- 0.0709100216627121
	pesos_i(6745) := b"0000000000000000_0000000000000000_0011000110100111_1011010110000000"; -- 0.19396528601646423
	pesos_i(6746) := b"1111111111111111_1111111111111111_1110100011110110_0111000010100000"; -- -0.08998962491750717
	pesos_i(6747) := b"1111111111111111_1111111111111111_1100010000010101_1110110111000000"; -- -0.23404039442539215
	pesos_i(6748) := b"1111111111111111_1111111111111111_0111000001000011_1001011000000000"; -- -0.5614687204360962
	pesos_i(6749) := b"1111111111111111_1111111111111111_1110111110001111_1101111101000000"; -- -0.0642109364271164
	pesos_i(6750) := b"0000000000000000_0000000000000000_0011110000101101_0001001110000000"; -- 0.23506280779838562
	pesos_i(6751) := b"1111111111111111_1111111111111111_1010111000111001_0111001110000000"; -- -0.31943586468696594
	pesos_i(6752) := b"0000000000000000_0000000000000000_0010001111000111_0100011100000000"; -- 0.13975948095321655
	pesos_i(6753) := b"1111111111111111_1111111111111111_1101010010101001_1000100111000000"; -- -0.1692880541086197
	pesos_i(6754) := b"1111111111111111_1111111111111111_1011101110000001_1100101110000000"; -- -0.2675507366657257
	pesos_i(6755) := b"0000000000000000_0000000000000000_0001010110111110_1001111100100000"; -- 0.08493990451097488
	pesos_i(6756) := b"0000000000000000_0000000000000000_0001010111110011_0110101111000000"; -- 0.08574555814266205
	pesos_i(6757) := b"0000000000000000_0000000000000000_1000011101110010_0000011000000000"; -- 0.5290836095809937
	pesos_i(6758) := b"0000000000000000_0000000000000000_0011100100000000_1111110000000000"; -- 0.2226712703704834
	pesos_i(6759) := b"1111111111111111_1111111111111111_1100001100110000_0100001011000000"; -- -0.23754484951496124
	pesos_i(6760) := b"1111111111111111_1111111111111111_1111110110111110_1001000001001000"; -- -0.008810980245471
	pesos_i(6761) := b"0000000000000000_0000000000000000_0000001001110010_1010111010110100"; -- 0.009562415070831776
	pesos_i(6762) := b"0000000000000000_0000000000000000_0100110111000010_1101111110000000"; -- 0.3037547767162323
	pesos_i(6763) := b"0000000000000000_0000000000000000_0011001000001110_0010011010000000"; -- 0.19552841782569885
	pesos_i(6764) := b"0000000000000000_0000000000000000_0001001011011101_1110101111000000"; -- 0.0736987441778183
	pesos_i(6765) := b"1111111111111111_1111111111111111_1111011010011001_1111110001000000"; -- -0.03671287000179291
	pesos_i(6766) := b"1111111111111111_1111111111111111_1100000001111101_1111101101000000"; -- -0.24807767570018768
	pesos_i(6767) := b"0000000000000000_0000000000000000_0010101010110000_0000100001000000"; -- 0.1667485386133194
	pesos_i(6768) := b"0000000000000000_0000000000000000_0111000111100111_0111111100000000"; -- 0.444938600063324
	pesos_i(6769) := b"1111111111111111_1111111111111111_0111111100010101_1010001000000000"; -- -0.5035761594772339
	pesos_i(6770) := b"0000000000000000_0000000000000000_0000001001000101_0101100010000100"; -- 0.008870632387697697
	pesos_i(6771) := b"1111111111111111_1111111111111111_1000000101010101_1010001010000000"; -- -0.4947870671749115
	pesos_i(6772) := b"0000000000000000_0000000000000000_0000110110111111_0011011101110000"; -- 0.053698983043432236
	pesos_i(6773) := b"1111111111111111_1111111111111111_1100110111011101_0010110110000000"; -- -0.19584384560585022
	pesos_i(6774) := b"1111111111111111_1111111111111111_1000110011111101_0001011110000000"; -- -0.4492631256580353
	pesos_i(6775) := b"1111111111111111_1111111111111111_1111010110101110_0011101011110000"; -- -0.04031020775437355
	pesos_i(6776) := b"1111111111111111_1111111111111111_1100000101001010_1100000001000000"; -- -0.24495314061641693
	pesos_i(6777) := b"1111111111111111_1111111111111111_1110101111101000_0111011101000000"; -- -0.07848410308361053
	pesos_i(6778) := b"0000000000000000_0000000000000000_0001111011010101_0011000000000000"; -- 0.12044048309326172
	pesos_i(6779) := b"1111111111111111_1111111111111111_1110101001001100_1101110000000000"; -- -0.08476471900939941
	pesos_i(6780) := b"0000000000000000_0000000000000000_1000001010110011_0011111000000000"; -- 0.5105475187301636
	pesos_i(6781) := b"1111111111111111_1111111111111111_1111111010011001_1100111101001110"; -- -0.005465548951178789
	pesos_i(6782) := b"1111111111111111_1111111111111111_1101100011001101_0011101101000000"; -- -0.15311841666698456
	pesos_i(6783) := b"1111111111111111_1111111111111111_1100000100001000_0101100111000000"; -- -0.2459663301706314
	pesos_i(6784) := b"1111111111111111_1111111111111111_1110011110011100_1111011110100000"; -- -0.0952611193060875
	pesos_i(6785) := b"1111111111111111_1111111111111111_1111111001010010_1101011011000000"; -- -0.006548479199409485
	pesos_i(6786) := b"0000000000000000_0000000000000000_0010000010101110_1111011011000000"; -- 0.12766973674297333
	pesos_i(6787) := b"1111111111111111_1111111111111111_1110100110111111_1110010110000000"; -- -0.08691564202308655
	pesos_i(6788) := b"0000000000000000_0000000000000000_0000000111101001_1001001110111000"; -- 0.007470352575182915
	pesos_i(6789) := b"1111111111111111_1111111111111111_1111111010010100_0000001000001110"; -- -0.005554076749831438
	pesos_i(6790) := b"0000000000000000_0000000000000000_0100010111010101_0010101000000000"; -- 0.27278387546539307
	pesos_i(6791) := b"1111111111111111_1111111111111111_1011100001010100_0101110010000000"; -- -0.2799627482891083
	pesos_i(6792) := b"1111111111111111_1111111111111111_1111010111001111_1101100010000000"; -- -0.03979727625846863
	pesos_i(6793) := b"1111111111111111_1111111111111111_1111101101100100_0110011100111000"; -- -0.01799921877682209
	pesos_i(6794) := b"1111111111111111_1111111111111111_1101101101101110_0101010000000000"; -- -0.14284777641296387
	pesos_i(6795) := b"1111111111111111_1111111111111111_1101010101011010_0111101111000000"; -- -0.16658808290958405
	pesos_i(6796) := b"0000000000000000_0000000000000000_0011010000111010_1100001011000000"; -- 0.204021617770195
	pesos_i(6797) := b"1111111111111111_1111111111111111_1110100011011100_1010111000100000"; -- -0.09038268774747849
	pesos_i(6798) := b"0000000000000000_0000000000000000_0010000010110100_0110000001000000"; -- 0.12775231897830963
	pesos_i(6799) := b"1111111111111111_1111111111111111_1111110101111011_1110010101101000"; -- -0.009828245267271996
	pesos_i(6800) := b"0000000000000000_0000000000000000_0010100000011011_0010011101000000"; -- 0.15666432678699493
	pesos_i(6801) := b"0000000000000000_0000000000000000_0101111010110001_1000011000000000"; -- 0.3698962926864624
	pesos_i(6802) := b"0000000000000000_0000000000000000_0010000000100011_1111011100000000"; -- 0.12554877996444702
	pesos_i(6803) := b"1111111111111111_1111111111111111_1010111001000110_0110000100000000"; -- -0.3192386031150818
	pesos_i(6804) := b"0000000000000000_0000000000000000_0001100110001110_1101010011000000"; -- 0.09983567893505096
	pesos_i(6805) := b"0000000000000000_0000000000000000_0100010000000010_0011111000000000"; -- 0.2656592130661011
	pesos_i(6806) := b"1111111111111111_1111111111111111_1111111100000010_0111011111111110"; -- -0.0038685803301632404
	pesos_i(6807) := b"0000000000000000_0000000000000000_0010010101010110_0110010111000000"; -- 0.1458495706319809
	pesos_i(6808) := b"0000000000000000_0000000000000000_0010011110000101_1111011100000000"; -- 0.15438789129257202
	pesos_i(6809) := b"1111111111111111_1111111111111111_1110101101101000_0110100000100000"; -- -0.08043812960386276
	pesos_i(6810) := b"0000000000000000_0000000000000000_0011001010010011_0101101100000000"; -- 0.19756096601486206
	pesos_i(6811) := b"1111111111111111_1111111111111111_1010000111101000_1010110000000000"; -- -0.36754345893859863
	pesos_i(6812) := b"1111111111111111_1111111111111111_1111100100110110_1000010001101000"; -- -0.02651188336312771
	pesos_i(6813) := b"1111111111111111_1111111111111111_1100111101001010_0001010001000000"; -- -0.1902758926153183
	pesos_i(6814) := b"1111111111111111_1111111111111111_1101110010101101_0000111010000000"; -- -0.13798436522483826
	pesos_i(6815) := b"1111111111111111_1111111111111111_1011011100111111_0100110000000000"; -- -0.28419041633605957
	pesos_i(6816) := b"0000000000000000_0000000000000000_0001001000000001_1001010111100000"; -- 0.07033669203519821
	pesos_i(6817) := b"0000000000000000_0000000000000000_0110010111100000_1010000110000000"; -- 0.3979588449001312
	pesos_i(6818) := b"1111111111111111_1111111111111111_1100111100001011_0111110100000000"; -- -0.19123095273971558
	pesos_i(6819) := b"1111111111111111_1111111111111111_1101110000100110_1101000001000000"; -- -0.14003275334835052
	pesos_i(6820) := b"1111111111111111_1111111111111111_1100101001110111_0101111111000000"; -- -0.20911599695682526
	pesos_i(6821) := b"0000000000000000_0000000000000000_0011111000100111_0101101010000000"; -- 0.24278798699378967
	pesos_i(6822) := b"1111111111111111_1111111111111111_1101110101110111_0001110101000000"; -- -0.13490121066570282
	pesos_i(6823) := b"0000000000000000_0000000000000000_0000111010111001_0000110110100000"; -- 0.057511188089847565
	pesos_i(6824) := b"1111111111111111_1111111111111111_1111100011111001_1111000010010000"; -- -0.02743622288107872
	pesos_i(6825) := b"1111111111111111_1111111111111111_1001110100010000_1000110010000000"; -- -0.38646623492240906
	pesos_i(6826) := b"1111111111111111_1111111111111111_1111111000101010_0001001010100000"; -- -0.007170520722866058
	pesos_i(6827) := b"0000000000000000_0000000000000000_0000110011011100_1100100100110000"; -- 0.05024392530322075
	pesos_i(6828) := b"0000000000000000_0000000000000000_0000010001111100_1000111011110000"; -- 0.017525609582662582
	pesos_i(6829) := b"0000000000000000_0000000000000000_0000111111101100_1100010111110000"; -- 0.06220662221312523
	pesos_i(6830) := b"1111111111111111_1111111111111111_1101001000101101_1111011010000000"; -- -0.17898616194725037
	pesos_i(6831) := b"1111111111111111_1111111111111111_1111111000010101_0101010000011110"; -- -0.007487051654607058
	pesos_i(6832) := b"0000000000000000_0000000000000000_0010010011011011_1001000010000000"; -- 0.14397528767585754
	pesos_i(6833) := b"1111111111111111_1111111111111111_1111011101100100_0100010011000000"; -- -0.03362627327442169
	pesos_i(6834) := b"1111111111111111_1111111111111111_1111101101111110_1111100100101000"; -- -0.01759379170835018
	pesos_i(6835) := b"1111111111111111_1111111111111111_1011001010110110_0100101000000000"; -- -0.3019059896469116
	pesos_i(6836) := b"1111111111111111_1111111111111111_1101110011101011_1101101100000000"; -- -0.1370261311531067
	pesos_i(6837) := b"0000000000000000_0000000000000000_0001101011011010_1010010001100000"; -- 0.10489871352910995
	pesos_i(6838) := b"0000000000000000_0000000000000000_0101000011101011_0000000010000000"; -- 0.3160858452320099
	pesos_i(6839) := b"1111111111111111_1111111111111111_1010101111110011_0000111000000000"; -- -0.32832252979278564
	pesos_i(6840) := b"0000000000000000_0000000000000000_0000100010110001_0110111011100000"; -- 0.03395741432905197
	pesos_i(6841) := b"0000000000000000_0000000000000000_0000100011100011_0000110011010000"; -- 0.034714508801698685
	pesos_i(6842) := b"1111111111111111_1111111111111111_1111001000101011_1010111011110000"; -- -0.054020944982767105
	pesos_i(6843) := b"0000000000000000_0000000000000000_0000101010110101_1101010010100000"; -- 0.04183701425790787
	pesos_i(6844) := b"1111111111111111_1111111111111111_1111000110000100_1100100111000000"; -- -0.056567564606666565
	pesos_i(6845) := b"0000000000000000_0000000000000000_0101000110010110_1111011010000000"; -- 0.31870976090431213
	pesos_i(6846) := b"1111111111111111_1111111111111111_1111000100111011_0010110111110000"; -- -0.05769074335694313
	pesos_i(6847) := b"1111111111111111_1111111111111111_1100111111001010_0010111101000000"; -- -0.18832115828990936
	pesos_i(6848) := b"1111111111111111_1111111111111111_1101101101001000_1010001100000000"; -- -0.1434229016304016
	pesos_i(6849) := b"1111111111111111_1111111111111111_1001101011011101_0111110000000000"; -- -0.39505791664123535
	pesos_i(6850) := b"0000000000000000_0000000000000000_0010000010011110_0001000001000000"; -- 0.1274118572473526
	pesos_i(6851) := b"0000000000000000_0000000000000000_0011010011001111_1111111111000000"; -- 0.2062988132238388
	pesos_i(6852) := b"1111111111111111_1111111111111111_1110010000001001_0011000100000000"; -- -0.1092347502708435
	pesos_i(6853) := b"0000000000000000_0000000000000000_0001110100101000_0000111011000000"; -- 0.11389248073101044
	pesos_i(6854) := b"1111111111111111_1111111111111111_0001001010001000_0110110100000000"; -- -0.9276058077812195
	pesos_i(6855) := b"0000000000000000_0000000000000000_0011001111101011_0110111101000000"; -- 0.20281119644641876
	pesos_i(6856) := b"0000000000000000_0000000000000000_0010111010100111_0000001100000000"; -- 0.18223589658737183
	pesos_i(6857) := b"0000000000000000_0000000000000000_0010110010100100_0011011111000000"; -- 0.17438076436519623
	pesos_i(6858) := b"1111111111111111_1111111111111111_1111000111001111_0110100111110000"; -- -0.05542886629700661
	pesos_i(6859) := b"0000000000000000_0000000000000000_0001010110101001_0101101100100000"; -- 0.08461541682481766
	pesos_i(6860) := b"0000000000000000_0000000000000000_0011110111101000_1011011110000000"; -- 0.24183222651481628
	pesos_i(6861) := b"1111111111111111_1111111111111111_1111111110110111_0011101101111100"; -- -0.0011103461729362607
	pesos_i(6862) := b"0000000000000000_0000000000000000_0100101110001111_1110001100000000"; -- 0.2951642870903015
	pesos_i(6863) := b"1111111111111111_1111111111111111_1101100011010000_0010010101000000"; -- -0.15307395160198212
	pesos_i(6864) := b"1111111111111111_1111111111111111_1101001110110100_1101011000000000"; -- -0.17302191257476807
	pesos_i(6865) := b"0000000000000000_0000000000000000_0001100011111011_1111010000000000"; -- 0.0975944995880127
	pesos_i(6866) := b"0000000000000000_0000000000000000_0100011000011100_1101101010000000"; -- 0.2738777697086334
	pesos_i(6867) := b"0000000000000000_0000000000000000_0000010011001110_1100111100111000"; -- 0.01878066174685955
	pesos_i(6868) := b"1111111111111111_1111111111111111_1101101000001001_0010110000000000"; -- -0.14829754829406738
	pesos_i(6869) := b"0000000000000000_0000000000000000_0001010010011111_0111110010100000"; -- 0.08055857568979263
	pesos_i(6870) := b"1111111111111111_1111111111111111_1101010010110111_0011111010000000"; -- -0.16907891631126404
	pesos_i(6871) := b"0000000000000000_0000000000000000_0000110000001000_0100111111100000"; -- 0.047001831233501434
	pesos_i(6872) := b"1111111111111111_1111111111111111_1111100110100011_0101110100000000"; -- -0.02485102415084839
	pesos_i(6873) := b"1111111111111111_1111111111111111_1110110000011001_0101000000100000"; -- -0.07773875445127487
	pesos_i(6874) := b"1111111111111111_1111111111111111_1111001000111101_1010110001010000"; -- -0.05374644324183464
	pesos_i(6875) := b"1111111111111111_1111111111111111_0101101110000010_0011110100000000"; -- -0.6425439715385437
	pesos_i(6876) := b"1111111111111111_1111111111111111_0000011011010000_1001111100000000"; -- -0.9733791947364807
	pesos_i(6877) := b"0000000000000000_0000000000000000_0001101101010001_1001011111000000"; -- 0.10671375691890717
	pesos_i(6878) := b"1111111111111111_1111111111111111_1011101101011110_0000010110000000"; -- -0.26809659600257874
	pesos_i(6879) := b"1111111111111111_1111111111111111_1101110010100101_1101010111000000"; -- -0.13809455931186676
	pesos_i(6880) := b"0000000000000000_0000000000000000_0011110100111111_0000100010000000"; -- 0.2392430603504181
	pesos_i(6881) := b"1111111111111111_1111111111111111_1101001011101100_0100111001000000"; -- -0.17608176171779633
	pesos_i(6882) := b"1111111111111111_1111111111111111_0111010100101100_1001101100000000"; -- -0.5422881245613098
	pesos_i(6883) := b"1111111111111111_1111111111111111_1101100001111011_0000100010000000"; -- -0.1543726623058319
	pesos_i(6884) := b"1111111111111111_1111111111111111_1010110000100100_0000000000000000"; -- -0.32757568359375
	pesos_i(6885) := b"0000000000000000_0000000000000000_0101010111100111_0010011010000000"; -- 0.33555832505226135
	pesos_i(6886) := b"1111111111111111_1111111111111111_1111000100000111_1100010000010000"; -- -0.058475252240896225
	pesos_i(6887) := b"0000000000000000_0000000000000000_0010101111000011_1000110001000000"; -- 0.17095257341861725
	pesos_i(6888) := b"0000000000000000_0000000000000000_0100100010001110_0010000100000000"; -- 0.2834187150001526
	pesos_i(6889) := b"1111111111111111_1111111111111111_1111010110101110_0111110111100000"; -- -0.0403062179684639
	pesos_i(6890) := b"0000000000000000_0000000000000000_0001001000000000_1111111111100000"; -- 0.0703277513384819
	pesos_i(6891) := b"1111111111111111_1111111111111111_1111100001011010_0101100101110000"; -- -0.0298713780939579
	pesos_i(6892) := b"0000000000000000_0000000000000000_0001110111000010_1110011110100000"; -- 0.1162552610039711
	pesos_i(6893) := b"1111111111111111_1111111111111111_1100110010101011_1101111100000000"; -- -0.2005024552345276
	pesos_i(6894) := b"1111111111111111_1111111111111111_1010110000100001_1111011000000000"; -- -0.32760679721832275
	pesos_i(6895) := b"0000000000000000_0000000000000000_0011111001010111_0010010110000000"; -- 0.24351724982261658
	pesos_i(6896) := b"0000000000000000_0000000000000000_0011110001110101_0100010001000000"; -- 0.23616434633731842
	pesos_i(6897) := b"1111111111111111_1111111111111111_1000010011110010_1110100110000000"; -- -0.48066845536231995
	pesos_i(6898) := b"1111111111111111_1111111111111111_1110101110001011_1100001111000000"; -- -0.07989861071109772
	pesos_i(6899) := b"0000000000000000_0000000000000000_0001111010111100_0001111001100000"; -- 0.12005796283483505
	pesos_i(6900) := b"0000000000000000_0000000000000000_0000100000100101_1010100110000000"; -- 0.03182467818260193
	pesos_i(6901) := b"1111111111111111_1111111111111111_1110100110010100_1100010011100000"; -- -0.08757371455430984
	pesos_i(6902) := b"0000000000000000_0000000000000000_0010100010111110_0110011110000000"; -- 0.15915533900260925
	pesos_i(6903) := b"0000000000000000_0000000000000000_0010010110011011_1001001010000000"; -- 0.1469050943851471
	pesos_i(6904) := b"0000000000000000_0000000000000000_0001000110001000_1001001101000000"; -- 0.06849022209644318
	pesos_i(6905) := b"1111111111111111_1111111111111111_1010101000101001_1111010000000000"; -- -0.3352973461151123
	pesos_i(6906) := b"0000000000000000_0000000000000000_0000111100101011_0010111101010000"; -- 0.059252697974443436
	pesos_i(6907) := b"0000000000000000_0000000000000000_0011010010010011_0110000111000000"; -- 0.2053738683462143
	pesos_i(6908) := b"0000000000000000_0000000000000000_0011010000000110_0100111101000000"; -- 0.20322127640247345
	pesos_i(6909) := b"0000000000000000_0000000000000000_0001100111110100_0100111111000000"; -- 0.10138414800167084
	pesos_i(6910) := b"0000000000000000_0000000000000000_0010011101100101_0001000001000000"; -- 0.1538858562707901
	pesos_i(6911) := b"1111111111111111_1111111111111111_1101111110010100_0010101000000000"; -- -0.12664544582366943
	pesos_i(6912) := b"0000000000000000_0000000000000000_0000010000111000_0101000111001000"; -- 0.016484366729855537
	pesos_i(6913) := b"1111111111111111_1111111111111111_1110010011010010_0000110001000000"; -- -0.1061699241399765
	pesos_i(6914) := b"0000000000000000_0000000000000000_0001000110000101_0100111100000000"; -- 0.06844037771224976
	pesos_i(6915) := b"1111111111111111_1111111111111111_1111110010100111_1111101001101000"; -- -0.013061856850981712
	pesos_i(6916) := b"0000000000000000_0000000000000000_0000101001011100_1110011101010000"; -- 0.04048009589314461
	pesos_i(6917) := b"0000000000000000_0000000000000000_0010101000110011_0011010010000000"; -- 0.1648438274860382
	pesos_i(6918) := b"0000000000000000_0000000000000000_0011101110001101_0110011110000000"; -- 0.23262640833854675
	pesos_i(6919) := b"1111111111111111_1111111111111111_1110000010111011_0110001011100000"; -- -0.12214071303606033
	pesos_i(6920) := b"1111111111111111_1111111111111111_1110100010001101_1110110100000000"; -- -0.09158438444137573
	pesos_i(6921) := b"0000000000000000_0000000000000000_0101010110010101_0100001110000000"; -- 0.33430883288383484
	pesos_i(6922) := b"1111111111111111_1111111111111111_1101100111001110_0010100100000000"; -- -0.1491979956626892
	pesos_i(6923) := b"1111111111111111_1111111111111111_1000111110010110_1110000010000000"; -- -0.4391040503978729
	pesos_i(6924) := b"1111111111111111_1111111111111111_1111111110111111_0001100111111110"; -- -0.0009902720339596272
	pesos_i(6925) := b"0000000000000000_0000000000000000_0001111001011001_0111010101000000"; -- 0.11855252087116241
	pesos_i(6926) := b"0000000000000000_0000000000000000_0001100011101011_1000111110100000"; -- 0.09734437614679337
	pesos_i(6927) := b"1111111111111111_1111111111111111_1100001000110011_1101011100000000"; -- -0.2413964867591858
	pesos_i(6928) := b"0000000000000000_0000000000000000_0100000111010111_0000010000000000"; -- 0.2571871280670166
	pesos_i(6929) := b"0000000000000000_0000000000000000_0010001010110000_0000111100000000"; -- 0.13549894094467163
	pesos_i(6930) := b"0000000000000000_0000000000000000_0000101010010010_1111100001100000"; -- 0.04130508750677109
	pesos_i(6931) := b"0000000000000000_0000000000000000_0010010001101000_1011001110000000"; -- 0.14222261309623718
	pesos_i(6932) := b"0000000000000000_0000000000000000_0001011110011100_1000101011000000"; -- 0.09223239123821259
	pesos_i(6933) := b"0000000000000000_0000000000000000_0000000010111110_1101101100110011"; -- 0.002912235213443637
	pesos_i(6934) := b"1111111111111111_1111111111111111_1111001001010010_0111011101010000"; -- -0.053429167717695236
	pesos_i(6935) := b"0000000000000000_0000000000000000_0001101000011010_1010101100100000"; -- 0.10196942836046219
	pesos_i(6936) := b"0000000000000000_0000000000000000_0001110110011101_1100110010100000"; -- 0.11568907648324966
	pesos_i(6937) := b"0000000000000000_0000000000000000_0010001101000001_1100111010000000"; -- 0.13772287964820862
	pesos_i(6938) := b"0000000000000000_0000000000000000_0011010001000011_1111010100000000"; -- 0.20416194200515747
	pesos_i(6939) := b"1111111111111111_1111111111111111_0110011101100000_1100110000000000"; -- -0.5961792469024658
	pesos_i(6940) := b"0000000000000000_0000000000000000_0001100011100101_1001011000000000"; -- 0.09725320339202881
	pesos_i(6941) := b"0000000000000000_0000000000000000_0001110111101100_0010111111000000"; -- 0.11688517034053802
	pesos_i(6942) := b"1111111111111111_1111111111111111_1101001111110011_1010010000000000"; -- -0.17206358909606934
	pesos_i(6943) := b"1111111111111111_1111111111111111_1010110011110101_0011111010000000"; -- -0.32438287138938904
	pesos_i(6944) := b"1111111111111111_1111111111111111_1011100011011001_0011000000000000"; -- -0.2779359817504883
	pesos_i(6945) := b"0000000000000000_0000000000000000_0011101010101110_0011010110000000"; -- 0.22922071814537048
	pesos_i(6946) := b"1111111111111111_1111111111111111_1010101110101100_1101101110000000"; -- -0.3293936550617218
	pesos_i(6947) := b"1111111111111111_1111111111111111_1110111110101101_0000110001100000"; -- -0.0637657418847084
	pesos_i(6948) := b"1111111111111111_1111111111111111_1101011001100110_0101110000000000"; -- -0.16250061988830566
	pesos_i(6949) := b"0000000000000000_0000000000000000_0001011111001001_1000110000000000"; -- 0.09291911125183105
	pesos_i(6950) := b"1111111111111111_1111111111111111_1010010110101000_1101110010000000"; -- -0.352892130613327
	pesos_i(6951) := b"0000000000000000_0000000000000000_0011010101011101_0100000111000000"; -- 0.20845423638820648
	pesos_i(6952) := b"0000000000000000_0000000000000000_0010000101101010_0011011101000000"; -- 0.13052697479724884
	pesos_i(6953) := b"1111111111111111_1111111111111111_1110001001001110_1111101001100000"; -- -0.11598239094018936
	pesos_i(6954) := b"1111111111111111_1111111111111111_1010001101001111_1010001010000000"; -- -0.3620661199092865
	pesos_i(6955) := b"1111111111111111_1111111111111111_1110111100110000_1100011100100000"; -- -0.0656619593501091
	pesos_i(6956) := b"1111111111111111_1111111111111111_1110111111111001_1010100011000000"; -- -0.06259675323963165
	pesos_i(6957) := b"1111111111111111_1111111111111111_1111111000101110_0110100100101110"; -- -0.007104326505213976
	pesos_i(6958) := b"1111111111111111_1111111111111111_1110101100111100_0011010111100000"; -- -0.08111251145601273
	pesos_i(6959) := b"0000000000000000_0000000000000000_0000110001101010_1111011010110000"; -- 0.04850713536143303
	pesos_i(6960) := b"0000000000000000_0000000000000000_0000000100101100_1111010001001100"; -- 0.004592197947204113
	pesos_i(6961) := b"1111111111111111_1111111111111111_1010001100100100_1000101110000000"; -- -0.36272361874580383
	pesos_i(6962) := b"1111111111111111_1111111111111111_1100010111101010_1010010011000000"; -- -0.22688837349414825
	pesos_i(6963) := b"1111111111111111_1111111111111111_1111111010100100_1101101010010100"; -- -0.005297030322253704
	pesos_i(6964) := b"1111111111111111_1111111111111111_1101101011100000_0010110101000000"; -- -0.1450168341398239
	pesos_i(6965) := b"1111111111111111_1111111111111111_1101011010100001_0100101000000000"; -- -0.16160142421722412
	pesos_i(6966) := b"0000000000000000_0000000000000000_0001110010101101_0010011000000000"; -- 0.11201703548431396
	pesos_i(6967) := b"1111111111111111_1111111111111111_1011010100010000_0010011000000000"; -- -0.29272234439849854
	pesos_i(6968) := b"0000000000000000_0000000000000000_0000101010101001_1101000100000000"; -- 0.04165369272232056
	pesos_i(6969) := b"0000000000000000_0000000000000000_0001100000101011_1011101010000000"; -- 0.09441724419593811
	pesos_i(6970) := b"0000000000000000_0000000000000000_0001010001111110_0100011000000000"; -- 0.08005177974700928
	pesos_i(6971) := b"1111111111111111_1111111111111111_1001011110000110_1101111000000000"; -- -0.40809834003448486
	pesos_i(6972) := b"1111111111111111_1111111111111111_1101001111101000_0111010111000000"; -- -0.1722341924905777
	pesos_i(6973) := b"0000000000000000_0000000000000000_0010010110001110_1101111010000000"; -- 0.14671126008033752
	pesos_i(6974) := b"0000000000000000_0000000000000000_0000001111010110_1000010001110000"; -- 0.01499202474951744
	pesos_i(6975) := b"1111111111111111_1111111111111111_1110101010000111_1011111000100000"; -- -0.08386623114347458
	pesos_i(6976) := b"1111111111111111_1111111111111111_1111000001100100_0000100011110000"; -- -0.06097358837723732
	pesos_i(6977) := b"1111111111111111_1111111111111111_1110000000001001_0100001011000000"; -- -0.12485869228839874
	pesos_i(6978) := b"0000000000000000_0000000000000000_0101010100101110_1010101110000000"; -- 0.332743376493454
	pesos_i(6979) := b"0000000000000000_0000000000000000_0010100010010111_0101110100000000"; -- 0.1585596203804016
	pesos_i(6980) := b"1111111111111111_1111111111111111_1010110001100100_1000001110000000"; -- -0.32659128308296204
	pesos_i(6981) := b"0000000000000000_0000000000000000_0000010011100110_1100101100111000"; -- 0.01914663426578045
	pesos_i(6982) := b"1111111111111111_1111111111111111_1011110010011011_0010111110000000"; -- -0.26325705647468567
	pesos_i(6983) := b"1111111111111111_1111111111111111_1101010001001110_0001001100000000"; -- -0.17068368196487427
	pesos_i(6984) := b"0000000000000000_0000000000000000_0001110100000111_1011001010100000"; -- 0.1133987084031105
	pesos_i(6985) := b"0000000000000000_0000000000000000_0011110010100100_1000001110000000"; -- 0.23688527941703796
	pesos_i(6986) := b"0000000000000000_0000000000000000_0001000111000111_0010001111100000"; -- 0.06944488734006882
	pesos_i(6987) := b"1111111111111111_1111111111111111_1100001011100110_1010101010000000"; -- -0.2386678159236908
	pesos_i(6988) := b"0000000000000000_0000000000000000_0010011000011101_1000010110000000"; -- 0.14888796210289001
	pesos_i(6989) := b"1111111111111111_1111111111111111_1111010001011000_1001110010010000"; -- -0.04552289471030235
	pesos_i(6990) := b"1111111111111111_1111111111111111_1110000111111101_0101000011100000"; -- -0.11722845584154129
	pesos_i(6991) := b"1111111111111111_1111111111111111_1110001101111110_0101101011100000"; -- -0.11135322600603104
	pesos_i(6992) := b"0000000000000000_0000000000000000_0001101110001110_1101000010000000"; -- 0.10764792561531067
	pesos_i(6993) := b"0000000000000000_0000000000000000_0100001100010011_1100110000000000"; -- 0.2620208263397217
	pesos_i(6994) := b"0000000000000000_0000000000000000_0011111100111011_1111110000000000"; -- 0.2470090389251709
	pesos_i(6995) := b"0000000000000000_0000000000000000_0101001110010001_0110011110000000"; -- 0.32643744349479675
	pesos_i(6996) := b"1111111111111111_1111111111111111_1101101101110001_1101111110000000"; -- -0.1427936851978302
	pesos_i(6997) := b"0000000000000000_0000000000000000_0001011000001110_0101101100000000"; -- 0.08615654706954956
	pesos_i(6998) := b"1111111111111111_1111111111111111_1100010011110000_1101100011000000"; -- -0.23069997131824493
	pesos_i(6999) := b"0000000000000000_0000000000000000_0011010100111011_1100100100000000"; -- 0.20794349908828735
	pesos_i(7000) := b"1111111111111111_1111111111111111_1100001100000100_1000110101000000"; -- -0.23821179568767548
	pesos_i(7001) := b"1111111111111111_1111111111111111_1011111110111100_1001001000000000"; -- -0.2510288953781128
	pesos_i(7002) := b"1111111111111111_1111111111111111_1100111001010110_1111000100000000"; -- -0.19398587942123413
	pesos_i(7003) := b"1111111111111111_1111111111111111_1111010001110101_1110001000010000"; -- -0.04507624730467796
	pesos_i(7004) := b"1111111111111111_1111111111111111_1000000011001101_1000000010000000"; -- -0.49686428904533386
	pesos_i(7005) := b"0000000000000000_0000000000000000_0000110111101000_0100101110100000"; -- 0.05432579666376114
	pesos_i(7006) := b"1111111111111111_1111111111111111_1010110110101001_1111100110000000"; -- -0.32162514328956604
	pesos_i(7007) := b"1111111111111111_1111111111111111_1111000011000001_0010000100100000"; -- -0.059553079307079315
	pesos_i(7008) := b"0000000000000000_0000000000000000_0100010111001101_0011110110000000"; -- 0.2726629674434662
	pesos_i(7009) := b"0000000000000000_0000000000000000_0001111001001111_0011001101000000"; -- 0.11839599907398224
	pesos_i(7010) := b"1111111111111111_1111111111111111_1000100011010110_1100101110000000"; -- -0.4654724895954132
	pesos_i(7011) := b"0000000000000000_0000000000000000_0000000111111011_1010010010001010"; -- 0.007746013347059488
	pesos_i(7012) := b"1111111111111111_1111111111111111_1101100110100110_0000010111000000"; -- -0.14981044828891754
	pesos_i(7013) := b"0000000000000000_0000000000000000_0010011111110001_0001011000000000"; -- 0.15602242946624756
	pesos_i(7014) := b"1111111111111111_1111111111111111_1110001110000111_1110100000000000"; -- -0.11120748519897461
	pesos_i(7015) := b"0000000000000000_0000000000000000_0001110011100110_1110100011000000"; -- 0.11289839446544647
	pesos_i(7016) := b"0000000000000000_0000000000000000_0011001001110001_1110001000000000"; -- 0.19705021381378174
	pesos_i(7017) := b"1111111111111111_1111111111111111_1110111110000001_0001010000000000"; -- -0.06443667411804199
	pesos_i(7018) := b"0000000000000000_0000000000000000_0001010110110010_0001000110000000"; -- 0.08474835753440857
	pesos_i(7019) := b"1111111111111111_1111111111111111_1111011010011001_1101010111110000"; -- -0.036715153604745865
	pesos_i(7020) := b"1111111111111111_1111111111111111_1111000001001100_0000111000110000"; -- -0.06133948639035225
	pesos_i(7021) := b"1111111111111111_1111111111111111_1110101101001000_0000100010100000"; -- -0.08093210309743881
	pesos_i(7022) := b"0000000000000000_0000000000000000_0000101001110010_0010011011000000"; -- 0.040804311633110046
	pesos_i(7023) := b"0000000000000000_0000000000000000_0001000000101010_0101000100000000"; -- 0.0631456971168518
	pesos_i(7024) := b"0000000000000000_0000000000000000_0100010010000111_0100101110000000"; -- 0.26768943667411804
	pesos_i(7025) := b"1111111111111111_1111111111111111_1101011111101100_0011110011000000"; -- -0.1565515547990799
	pesos_i(7026) := b"0000000000000000_0000000000000000_0001000111100110_1111010011000000"; -- 0.06993035972118378
	pesos_i(7027) := b"1111111111111111_1111111111111111_1100101100011000_0101011001000000"; -- -0.20665989816188812
	pesos_i(7028) := b"0000000000000000_0000000000000000_0010111000101110_0111111010000000"; -- 0.1803969442844391
	pesos_i(7029) := b"1111111111111111_1111111111111111_1100111010111110_1100101011000000"; -- -0.1924012452363968
	pesos_i(7030) := b"0000000000000000_0000000000000000_0001000000101111_0000100101100000"; -- 0.06321772187948227
	pesos_i(7031) := b"0000000000000000_0000000000000000_0001001010111110_0110110111000000"; -- 0.0732182115316391
	pesos_i(7032) := b"0000000000000000_0000000000000000_0000100100011110_1100100111100000"; -- 0.03562604635953903
	pesos_i(7033) := b"1111111111111111_1111111111111111_1000101110010100_1101100000000000"; -- -0.4547600746154785
	pesos_i(7034) := b"0000000000000000_0000000000000000_0001100000011010_0010110100000000"; -- 0.09414941072463989
	pesos_i(7035) := b"1111111111111111_1111111111111111_1110011001000101_1110011111000000"; -- -0.1004958301782608
	pesos_i(7036) := b"1111111111111111_1111111111111111_1111110000100110_1100010011010100"; -- -0.015033434145152569
	pesos_i(7037) := b"1111111111111111_1111111111111111_1111011110110111_0000001100100000"; -- -0.03236370533704758
	pesos_i(7038) := b"0000000000000000_0000000000000000_0011011001000000_0001101111000000"; -- 0.21191571652889252
	pesos_i(7039) := b"0000000000000000_0000000000000000_0011001000000101_0100101111000000"; -- 0.19539330899715424
	pesos_i(7040) := b"0000000000000000_0000000000000000_0000010110101101_0101001001101000"; -- 0.022175932303071022
	pesos_i(7041) := b"0000000000000000_0000000000000000_0011100010100010_1011111100000000"; -- 0.2212333083152771
	pesos_i(7042) := b"0000000000000000_0000000000000000_0010100010101001_1001000110000000"; -- 0.15883740782737732
	pesos_i(7043) := b"0000000000000000_0000000000000000_0010010111110000_1101001001000000"; -- 0.14820589125156403
	pesos_i(7044) := b"0000000000000000_0000000000000000_0001010001100011_0001101101100000"; -- 0.07963725179433823
	pesos_i(7045) := b"1111111111111111_1111111111111111_1111010001101110_1100000001110000"; -- -0.045185063034296036
	pesos_i(7046) := b"0000000000000000_0000000000000000_0001001000100111_1111100001000000"; -- 0.07092238962650299
	pesos_i(7047) := b"0000000000000000_0000000000000000_0001110001111011_1100011011000000"; -- 0.11126367747783661
	pesos_i(7048) := b"0000000000000000_0000000000000000_0000110100001010_1010000101100000"; -- 0.05094345659017563
	pesos_i(7049) := b"0000000000000000_0000000000000000_0011110110101000_0110110010000000"; -- 0.24085119366645813
	pesos_i(7050) := b"1111111111111111_1111111111111111_1011111111011010_0011111100000000"; -- -0.25057607889175415
	pesos_i(7051) := b"1111111111111111_1111111111111111_1100100111011100_0011010010000000"; -- -0.2114836871623993
	pesos_i(7052) := b"1111111111111111_1111111111111111_1101111110001001_0111100111000000"; -- -0.1268085390329361
	pesos_i(7053) := b"1111111111111111_1111111111111111_1110000010100010_1111111011000000"; -- -0.12251289188861847
	pesos_i(7054) := b"1111111111111111_1111111111111111_1101100101111110_0001100110000000"; -- -0.15041962265968323
	pesos_i(7055) := b"1111111111111111_1111111111111111_1111110111000100_0011100010100100"; -- -0.008724651299417019
	pesos_i(7056) := b"0000000000000000_0000000000000000_0010011000110110_1101100000000000"; -- 0.14927434921264648
	pesos_i(7057) := b"0000000000000000_0000000000000000_0000101010111011_1100001001100000"; -- 0.04192747920751572
	pesos_i(7058) := b"0000000000000000_0000000000000000_0100111110100010_1011110100000000"; -- 0.31107693910598755
	pesos_i(7059) := b"0000000000000000_0000000000000000_0000001001001110_1110110111000100"; -- 0.009016857482492924
	pesos_i(7060) := b"0000000000000000_0000000000000000_0000010000000101_1010011011000000"; -- 0.015711233019828796
	pesos_i(7061) := b"0000000000000000_0000000000000000_0001001001110000_0000100001100000"; -- 0.0720219835639
	pesos_i(7062) := b"0000000000000000_0000000000000000_0000001100000011_1010000101010000"; -- 0.01177414134144783
	pesos_i(7063) := b"0000000000000000_0000000000000000_0011000101100100_0111001001000000"; -- 0.1929389387369156
	pesos_i(7064) := b"0000000000000000_0000000000000000_0001000001011101_0100001000100000"; -- 0.06392300873994827
	pesos_i(7065) := b"1111111111111111_1111111111111111_1110110010110001_1011010010000000"; -- -0.07541343569755554
	pesos_i(7066) := b"0000000000000000_0000000000000000_0000101010100011_0100010000000000"; -- 0.04155373573303223
	pesos_i(7067) := b"1111111111111111_1111111111111111_1110111111000000_0100011001000000"; -- -0.06347237527370453
	pesos_i(7068) := b"1111111111111111_1111111111111111_1101100010001111_0011011110000000"; -- -0.15406468510627747
	pesos_i(7069) := b"1111111111111111_1111111111111111_1111010011011010_1100001011100000"; -- -0.043536968529224396
	pesos_i(7070) := b"0000000000000000_0000000000000000_0000001100010100_0101101111101100"; -- 0.012029404751956463
	pesos_i(7071) := b"1111111111111111_1111111111111111_1111101111110110_0011110010000000"; -- -0.01577398180961609
	pesos_i(7072) := b"1111111111111111_1111111111111111_1010100100010111_1111100110000000"; -- -0.33947792649269104
	pesos_i(7073) := b"0000000000000000_0000000000000000_0011010110000011_0001001010000000"; -- 0.20903125405311584
	pesos_i(7074) := b"0000000000000000_0000000000000000_0000101011011110_1110101010000000"; -- 0.04246392846107483
	pesos_i(7075) := b"1111111111111111_1111111111111111_1110110101110011_0001010000100000"; -- -0.0724627897143364
	pesos_i(7076) := b"1111111111111111_1111111111111111_1111111111011001_0000111010111010"; -- -0.000594214943703264
	pesos_i(7077) := b"0000000000000000_0000000000000000_0000011010111010_0010011111100000"; -- 0.02627801150083542
	pesos_i(7078) := b"1111111111111111_1111111111111111_1111110101011000_0100000101111100"; -- -0.010372073389589787
	pesos_i(7079) := b"0000000000000000_0000000000000000_0001011100100000_0000100000100000"; -- 0.0903325155377388
	pesos_i(7080) := b"0000000000000000_0000000000000000_0010101110010001_0000111010000000"; -- 0.17018213868141174
	pesos_i(7081) := b"0000000000000000_0000000000000000_0010000111001110_1010100111000000"; -- 0.13205967843532562
	pesos_i(7082) := b"1111111111111111_1111111111111111_1011100101011100_0011010000000000"; -- -0.2759368419647217
	pesos_i(7083) := b"0000000000000000_0000000000000000_0011011111101101_0011001010000000"; -- 0.21846309304237366
	pesos_i(7084) := b"0000000000000000_0000000000000000_0010111001111011_0010110101000000"; -- 0.1815670281648636
	pesos_i(7085) := b"0000000000000000_0000000000000000_0001101010101100_0100110001000000"; -- 0.10419155657291412
	pesos_i(7086) := b"0000000000000000_0000000000000000_0010000010001011_0100110000000000"; -- 0.12712550163269043
	pesos_i(7087) := b"1111111111111111_1111111111111111_1111100010010100_0011001100001000"; -- -0.028988657519221306
	pesos_i(7088) := b"0000000000000000_0000000000000000_0000110111111111_0100111001000000"; -- 0.054676905274391174
	pesos_i(7089) := b"1111111111111111_1111111111111111_1111001011011000_1110100001000000"; -- -0.051377758383750916
	pesos_i(7090) := b"1111111111111111_1111111111111111_1110111110000000_0001111110100000"; -- -0.06445124000310898
	pesos_i(7091) := b"0000000000000000_0000000000000000_0001001100110110_0101010000100000"; -- 0.07504773885011673
	pesos_i(7092) := b"1111111111111111_1111111111111111_1111111110001001_1101011110110110"; -- -0.0018029386410489678
	pesos_i(7093) := b"1111111111111111_1111111111111111_1110110011110010_1011101110100000"; -- -0.07442118972539902
	pesos_i(7094) := b"1111111111111111_1111111111111111_1111011010001111_0010011101000000"; -- -0.036878153681755066
	pesos_i(7095) := b"1111111111111111_1111111111111111_1110110001011001_0101010110000000"; -- -0.0767618715763092
	pesos_i(7096) := b"1111111111111111_1111111111111111_1111000011101111_0110101111100000"; -- -0.058846719563007355
	pesos_i(7097) := b"0000000000000000_0000000000000000_0001111100000100_0000110110100000"; -- 0.12115559726953506
	pesos_i(7098) := b"0000000000000000_0000000000000000_0001001001111110_1001100111100000"; -- 0.07224427908658981
	pesos_i(7099) := b"1111111111111111_1111111111111111_1110010001001001_1001111000000000"; -- -0.10825169086456299
	pesos_i(7100) := b"1111111111111111_1111111111111111_1101111100100000_1100001111000000"; -- -0.12840630114078522
	pesos_i(7101) := b"0000000000000000_0000000000000000_0011110110000011_0111000111000000"; -- 0.2402869313955307
	pesos_i(7102) := b"1111111111111111_1111111111111111_1110000101111001_0111011001100000"; -- -0.11924038082361221
	pesos_i(7103) := b"1111111111111111_1111111111111111_1111110000011110_0011001010100000"; -- -0.015164218842983246
	pesos_i(7104) := b"0000000000000000_0000000000000000_0010100011110101_1100101111000000"; -- 0.16000054776668549
	pesos_i(7105) := b"0000000000000000_0000000000000000_0000111000000000_1001011101010000"; -- 0.054696518927812576
	pesos_i(7106) := b"0000000000000000_0000000000000000_0001110010111100_1000110010100000"; -- 0.11225203424692154
	pesos_i(7107) := b"0000000000000000_0000000000000000_0011101000111000_0111001110000000"; -- 0.22742387652397156
	pesos_i(7108) := b"1111111111111111_1111111111111111_1100110000111101_1101100001000000"; -- -0.20218132436275482
	pesos_i(7109) := b"1111111111111111_1111111111111111_1111100111011000_1100110001010000"; -- -0.024035673588514328
	pesos_i(7110) := b"0000000000000000_0000000000000000_0010011111111100_0001000111000000"; -- 0.15619002282619476
	pesos_i(7111) := b"1111111111111111_1111111111111111_1110111000011010_0110110000100000"; -- -0.06990932673215866
	pesos_i(7112) := b"0000000000000000_0000000000000000_0010110010101110_0010110101000000"; -- 0.1745327264070511
	pesos_i(7113) := b"0000000000000000_0000000000000000_0000110111010000_1111100111000000"; -- 0.053969964385032654
	pesos_i(7114) := b"1111111111111111_1111111111111111_1111001011101011_1101010110110000"; -- -0.05108894780278206
	pesos_i(7115) := b"1111111111111111_1111111111111111_1110000001011001_1000100101100000"; -- -0.12363377958536148
	pesos_i(7116) := b"1111111111111111_1111111111111111_1110101101001011_0000000111100000"; -- -0.08088672906160355
	pesos_i(7117) := b"1111111111111111_1111111111111111_1110000101101010_1010111111000000"; -- -0.11946584284305573
	pesos_i(7118) := b"1111111111111111_1111111111111111_1101101111100100_1111110011000000"; -- -0.14103718101978302
	pesos_i(7119) := b"1111111111111111_1111111111111111_1110001100100001_1011000100100000"; -- -0.11276715248823166
	pesos_i(7120) := b"0000000000000000_0000000000000000_0010000011000001_0001111010000000"; -- 0.12794676423072815
	pesos_i(7121) := b"0000000000000000_0000000000000000_0010100111010000_0110010100000000"; -- 0.16333609819412231
	pesos_i(7122) := b"0000000000000000_0000000000000000_0001101010001001_0101010001000000"; -- 0.10365797579288483
	pesos_i(7123) := b"0000000000000000_0000000000000000_0001011011110100_0111101101000000"; -- 0.08966799080371857
	pesos_i(7124) := b"0000000000000000_0000000000000000_0000111010101111_0111101010010000"; -- 0.057365093380212784
	pesos_i(7125) := b"1111111111111111_1111111111111111_1110010110011101_0000001000000000"; -- -0.10307300090789795
	pesos_i(7126) := b"1111111111111111_1111111111111111_1101110010011001_0101000001000000"; -- -0.13828562200069427
	pesos_i(7127) := b"0000000000000000_0000000000000000_0010001100010110_1101011101000000"; -- 0.1370672732591629
	pesos_i(7128) := b"0000000000000000_0000000000000000_0000101101000110_1011010101000000"; -- 0.04404766857624054
	pesos_i(7129) := b"1111111111111111_1111111111111111_1110111100011011_1100010010100000"; -- -0.06598254293203354
	pesos_i(7130) := b"1111111111111111_1111111111111111_1110011100000100_0110100001000000"; -- -0.09758900105953217
	pesos_i(7131) := b"1111111111111111_1111111111111111_1110010000010001_0110011111100000"; -- -0.10910940915346146
	pesos_i(7132) := b"1111111111111111_1111111111111111_1101101000101111_1000100011000000"; -- -0.14771218597888947
	pesos_i(7133) := b"0000000000000000_0000000000000000_0000111101001111_1001011110100000"; -- 0.05980823189020157
	pesos_i(7134) := b"1111111111111111_1111111111111111_1011110100111100_0010101100000000"; -- -0.26080065965652466
	pesos_i(7135) := b"1111111111111111_1111111111111111_1111110111010111_1010101000110000"; -- -0.008427966386079788
	pesos_i(7136) := b"0000000000000000_0000000000000000_0100011111110001_1110100000000000"; -- 0.2810349464416504
	pesos_i(7137) := b"1111111111111111_1111111111111111_1101111110111101_0100110011000000"; -- -0.126017764210701
	pesos_i(7138) := b"1111111111111111_1111111111111111_1100110100011100_1111110101000000"; -- -0.19877640902996063
	pesos_i(7139) := b"1111111111111111_1111111111111111_1101000010001111_0111101010000000"; -- -0.18531069159507751
	pesos_i(7140) := b"1111111111111111_1111111111111111_1100100000010010_1101000110000000"; -- -0.21846285462379456
	pesos_i(7141) := b"0000000000000000_0000000000000000_0001100101100010_1100011110000000"; -- 0.09916350245475769
	pesos_i(7142) := b"1111111111111111_1111111111111111_1101000111011001_1001110100000000"; -- -0.18027323484420776
	pesos_i(7143) := b"0000000000000000_0000000000000000_0001101001000001_0110001001000000"; -- 0.10256017744541168
	pesos_i(7144) := b"1111111111111111_1111111111111111_1111000000001001_1110110100100000"; -- -0.062348537147045135
	pesos_i(7145) := b"0000000000000000_0000000000000000_0000010101000011_1000100101111000"; -- 0.020561782643198967
	pesos_i(7146) := b"0000000000000000_0000000000000000_0010101110001011_1111010010000000"; -- 0.17010429501533508
	pesos_i(7147) := b"0000000000000000_0000000000000000_0010111100001001_1000000101000000"; -- 0.18373878300189972
	pesos_i(7148) := b"1111111111111111_1111111111111111_1110001000001000_0010000111100000"; -- -0.11706341058015823
	pesos_i(7149) := b"0000000000000000_0000000000000000_0011100001100000_1101111101000000"; -- 0.2202281504869461
	pesos_i(7150) := b"0000000000000000_0000000000000000_0011001010100011_1110010100000000"; -- 0.19781333208084106
	pesos_i(7151) := b"0000000000000000_0000000000000000_0001011100010001_0001011000100000"; -- 0.09010446816682816
	pesos_i(7152) := b"1111111111111111_1111111111111111_1110010010011110_0100001111000000"; -- -0.10696007311344147
	pesos_i(7153) := b"0000000000000000_0000000000000000_0010001011110000_1000101111000000"; -- 0.13648293912410736
	pesos_i(7154) := b"1111111111111111_1111111111111111_1100011101111011_0000101000000000"; -- -0.22077882289886475
	pesos_i(7155) := b"0000000000000000_0000000000000000_0000110111110110_1110011101010000"; -- 0.05454869940876961
	pesos_i(7156) := b"0000000000000000_0000000000000000_0010010110000110_0111101010000000"; -- 0.14658322930335999
	pesos_i(7157) := b"0000000000000000_0000000000000000_0010101000010110_1101101101000000"; -- 0.164411261677742
	pesos_i(7158) := b"0000000000000000_0000000000000000_0011001000110110_1001011101000000"; -- 0.19614548981189728
	pesos_i(7159) := b"1111111111111111_1111111111111111_1100111111001100_0000101110000000"; -- -0.18829277157783508
	pesos_i(7160) := b"1111111111111111_1111111111111111_1011111001100011_0010100000000000"; -- -0.2562994956970215
	pesos_i(7161) := b"1111111111111111_1111111111111111_1100110011100100_1000001111000000"; -- -0.19963814318180084
	pesos_i(7162) := b"1111111111111111_1111111111111111_1111101001101000_1111011101101000"; -- -0.02183583937585354
	pesos_i(7163) := b"0000000000000000_0000000000000000_0001101101010101_0111011100100000"; -- 0.10677284747362137
	pesos_i(7164) := b"0000000000000000_0000000000000000_0000110111100100_0011000010100000"; -- 0.0542631521821022
	pesos_i(7165) := b"0000000000000000_0000000000000000_0001000010100100_1111011010000000"; -- 0.06501713395118713
	pesos_i(7166) := b"1111111111111111_1111111111111111_1111101010001010_0000010000100000"; -- -0.0213315412402153
	pesos_i(7167) := b"0000000000000000_0000000000000000_0011110011000011_0101111101000000"; -- 0.23735614120960236
	pesos_i(7168) := b"0000000000000000_0000000000000000_0001010110001111_1111110100100000"; -- 0.08422834426164627
	pesos_i(7169) := b"0000000000000000_0000000000000000_0101100111011010_0111011100000000"; -- 0.35098975896835327
	pesos_i(7170) := b"1111111111111111_1111111111111111_1101111010011111_1111101110000000"; -- -0.1303713619709015
	pesos_i(7171) := b"1111111111111111_1111111111111111_1101011001100001_1100111001000000"; -- -0.16257010400295258
	pesos_i(7172) := b"1111111111111111_1111111111111111_1011111110011010_0000001000000000"; -- -0.25155627727508545
	pesos_i(7173) := b"1111111111111111_1111111111111111_1110001111110101_1011010110000000"; -- -0.10953202843666077
	pesos_i(7174) := b"1111111111111111_1111111111111111_1110010100101000_0100010100100000"; -- -0.1048542782664299
	pesos_i(7175) := b"1111111111111111_1111111111111111_1101110011101000_1011101100000000"; -- -0.137073814868927
	pesos_i(7176) := b"1111111111111111_1111111111111111_1101000001100000_1101000110000000"; -- -0.18602266907691956
	pesos_i(7177) := b"1111111111111111_1111111111111111_1100010000001100_1010011110000000"; -- -0.23418191075325012
	pesos_i(7178) := b"1111111111111111_1111111111111111_1111111000011110_0001100111010000"; -- -0.007353197783231735
	pesos_i(7179) := b"1111111111111111_1111111111111111_1111100000001100_1001110000100000"; -- -0.031057588756084442
	pesos_i(7180) := b"0000000000000000_0000000000000000_0001000101000000_1010110011000000"; -- 0.06739310920238495
	pesos_i(7181) := b"0000000000000000_0000000000000000_0001000010000100_0101110001100000"; -- 0.06451966613531113
	pesos_i(7182) := b"0000000000000000_0000000000000000_0000000001010111_1000101010100110"; -- 0.0013357787393033504
	pesos_i(7183) := b"0000000000000000_0000000000000000_0001000111101000_0110001111000000"; -- 0.06995223462581635
	pesos_i(7184) := b"1111111111111111_1111111111111111_1110100000001000_0011011000000000"; -- -0.09362471103668213
	pesos_i(7185) := b"1111111111111111_1111111111111111_1011011010000010_1111001010000000"; -- -0.28706440329551697
	pesos_i(7186) := b"1111111111111111_1111111111111111_1110001111111011_0011001101000000"; -- -0.10944823920726776
	pesos_i(7187) := b"1111111111111111_1111111111111111_1101110000000011_1111010000000000"; -- -0.1405646800994873
	pesos_i(7188) := b"1111111111111111_1111111111111111_1101010101100110_1101000110000000"; -- -0.16639986634254456
	pesos_i(7189) := b"0000000000000000_0000000000000000_0001001101100101_0111001000000000"; -- 0.0757666826248169
	pesos_i(7190) := b"0000000000000000_0000000000000000_0001011111110110_1101100011100000"; -- 0.09361033886671066
	pesos_i(7191) := b"0000000000000000_0000000000000000_0001111110101000_1101001000000000"; -- 0.12366974353790283
	pesos_i(7192) := b"0000000000000000_0000000000000000_0001100011100010_1000100010100000"; -- 0.09720662981271744
	pesos_i(7193) := b"0000000000000000_0000000000000000_0101110001111100_0100010110000000"; -- 0.3612712323665619
	pesos_i(7194) := b"1111111111111111_1111111111111111_1111110001100100_1111000010101100"; -- -0.014084775932133198
	pesos_i(7195) := b"0000000000000000_0000000000000000_0010101100010111_1010101111000000"; -- 0.16832993924617767
	pesos_i(7196) := b"1111111111111111_1111111111111111_1101001000111011_0011101110000000"; -- -0.17878368496894836
	pesos_i(7197) := b"1111111111111111_1111111111111111_1110010001111110_0100100011000000"; -- -0.10744805634021759
	pesos_i(7198) := b"0000000000000000_0000000000000000_0010011101101101_0101001010000000"; -- 0.15401187539100647
	pesos_i(7199) := b"0000000000000000_0000000000000000_0000000111111001_1110111001111000"; -- 0.007719902321696281
	pesos_i(7200) := b"1111111111111111_1111111111111111_1111111000010101_1110000111001100"; -- -0.007478606887161732
	pesos_i(7201) := b"1111111111111111_1111111111111111_1111110101001010_1111101001100000"; -- -0.010574676096439362
	pesos_i(7202) := b"1111111111111111_1111111111111111_1110000101010011_1000001011100000"; -- -0.11981946974992752
	pesos_i(7203) := b"0000000000000000_0000000000000000_0011000011010110_0010011011000000"; -- 0.19076769053936005
	pesos_i(7204) := b"0000000000000000_0000000000000000_0000111110011111_0111101010100000"; -- 0.06102720648050308
	pesos_i(7205) := b"1111111111111111_1111111111111111_1011100101100001_0101010010000000"; -- -0.275858610868454
	pesos_i(7206) := b"1111111111111111_1111111111111111_1111011111101011_1000000110100000"; -- -0.03156270831823349
	pesos_i(7207) := b"0000000000000000_0000000000000000_0011100110010001_1000100000000000"; -- 0.22487688064575195
	pesos_i(7208) := b"0000000000000000_0000000000000000_0001000110011001_0011011110000000"; -- 0.06874415278434753
	pesos_i(7209) := b"1111111111111111_1111111111111111_1101000111111010_0010001010000000"; -- -0.17977699637413025
	pesos_i(7210) := b"0000000000000000_0000000000000000_0000001001001110_0111011111110000"; -- 0.009009834378957748
	pesos_i(7211) := b"0000000000000000_0000000000000000_0000100110110010_0111101101100000"; -- 0.037879668176174164
	pesos_i(7212) := b"0000000000000000_0000000000000000_0010010011111000_0101001000000000"; -- 0.14441406726837158
	pesos_i(7213) := b"1111111111111111_1111111111111111_1011010000101101_0001011000000000"; -- -0.29618704319000244
	pesos_i(7214) := b"1111111111111111_1111111111111111_1111001010111100_0100011010100000"; -- -0.05181463807821274
	pesos_i(7215) := b"1111111111111111_1111111111111111_1111010110111000_0111010111000000"; -- -0.0401541143655777
	pesos_i(7216) := b"1111111111111111_1111111111111111_1110000000001001_0110001011000000"; -- -0.12485678493976593
	pesos_i(7217) := b"1111111111111111_1111111111111111_1111011001101111_0010100010110000"; -- -0.0373663492500782
	pesos_i(7218) := b"1111111111111111_1111111111111111_1111000000001100_0101100100110000"; -- -0.062311578541994095
	pesos_i(7219) := b"0000000000000000_0000000000000000_0011001100001111_1111100011000000"; -- 0.19946245849132538
	pesos_i(7220) := b"0000000000000000_0000000000000000_0100001110001000_1010111110000000"; -- 0.2638044059276581
	pesos_i(7221) := b"0000000000000000_0000000000000000_0000101101101000_0110100010110000"; -- 0.044561903923749924
	pesos_i(7222) := b"1111111111111111_1111111111111111_1010100011101010_0111101010000000"; -- -0.34017214179039
	pesos_i(7223) := b"0000000000000000_0000000000000000_0011110000111111_0000110010000000"; -- 0.2353370487689972
	pesos_i(7224) := b"1111111111111111_1111111111111111_1101110100100110_1000000001000000"; -- -0.13613127171993256
	pesos_i(7225) := b"0000000000000000_0000000000000000_0001000101001110_0101110101000000"; -- 0.0676019936800003
	pesos_i(7226) := b"0000000000000000_0000000000000000_0100100010001010_1111100100000000"; -- 0.2833705544471741
	pesos_i(7227) := b"0000000000000000_0000000000000000_0001001111100000_0111000110000000"; -- 0.077643483877182
	pesos_i(7228) := b"0000000000000000_0000000000000000_0000110110011111_1110111101110000"; -- 0.05322166904807091
	pesos_i(7229) := b"1111111111111111_1111111111111111_1110100110110111_0011000011100000"; -- -0.0870484784245491
	pesos_i(7230) := b"0000000000000000_0000000000000000_0010000101111010_0011111110000000"; -- 0.13077160716056824
	pesos_i(7231) := b"1111111111111111_1111111111111111_1011100110010100_1010111100000000"; -- -0.2750750184059143
	pesos_i(7232) := b"1111111111111111_1111111111111111_1110010110000101_0001000011000000"; -- -0.10343833267688751
	pesos_i(7233) := b"0000000000000000_0000000000000000_0001100101101001_1000000001100000"; -- 0.09926607459783554
	pesos_i(7234) := b"1111111111111111_1111111111111111_1100001111001000_1001001000000000"; -- -0.2352207899093628
	pesos_i(7235) := b"1111111111111111_1111111111111111_1111011110010001_0010100010100000"; -- -0.0329413041472435
	pesos_i(7236) := b"1111111111111111_1111111111111111_1111000100000010_0110111101100000"; -- -0.05855659395456314
	pesos_i(7237) := b"0000000000000000_0000000000000000_0001000001000101_1000000101100000"; -- 0.06356056779623032
	pesos_i(7238) := b"1111111111111111_1111111111111111_1110100011001110_0100111101000000"; -- -0.09060196578502655
	pesos_i(7239) := b"1111111111111111_1111111111111111_1101011001000010_1001000000000000"; -- -0.16304683685302734
	pesos_i(7240) := b"1111111111111111_1111111111111111_1111011001111100_0010100111000000"; -- -0.03716792166233063
	pesos_i(7241) := b"0000000000000000_0000000000000000_0000001111011101_0010111110100000"; -- 0.015093781054019928
	pesos_i(7242) := b"0000000000000000_0000000000000000_0011011011100110_1001101101000000"; -- 0.21445627510547638
	pesos_i(7243) := b"0000000000000000_0000000000000000_0000001101111001_0111100001001000"; -- 0.01357223279774189
	pesos_i(7244) := b"1111111111111111_1111111111111111_1011001001101001_0001010100000000"; -- -0.3030840754508972
	pesos_i(7245) := b"0000000000000000_0000000000000000_0000101101101010_0111110110010000"; -- 0.04459366574883461
	pesos_i(7246) := b"1111111111111111_1111111111111111_1010110110011110_1100001000000000"; -- -0.3217962980270386
	pesos_i(7247) := b"1111111111111111_1111111111111111_1110000001001000_1000010101000000"; -- -0.12389342486858368
	pesos_i(7248) := b"0000000000000000_0000000000000000_0001111001011011_0010011101100000"; -- 0.11857839673757553
	pesos_i(7249) := b"0000000000000000_0000000000000000_0001000100000111_0111111110000000"; -- 0.06652066111564636
	pesos_i(7250) := b"1111111111111111_1111111111111111_1111001001000110_1000101011010000"; -- -0.053611110895872116
	pesos_i(7251) := b"1111111111111111_1111111111111111_1101000101110110_0010111101000000"; -- -0.18179039657115936
	pesos_i(7252) := b"0000000000000000_0000000000000000_0000000001001011_1001000010010110"; -- 0.0011530272895470262
	pesos_i(7253) := b"0000000000000000_0000000000000000_0100000001011101_0111010100000000"; -- 0.2514260411262512
	pesos_i(7254) := b"0000000000000000_0000000000000000_0101110010101000_1001010000000000"; -- 0.36194729804992676
	pesos_i(7255) := b"1111111111111111_1111111111111111_1101101111010010_0111101111000000"; -- -0.14131952822208405
	pesos_i(7256) := b"0000000000000000_0000000000000000_0010110100010101_0110101100000000"; -- 0.17610806226730347
	pesos_i(7257) := b"0000000000000000_0000000000000000_0000010000101001_0101101110101000"; -- 0.016256073489785194
	pesos_i(7258) := b"0000000000000000_0000000000000000_0000010111111011_1010010110101000"; -- 0.023371079936623573
	pesos_i(7259) := b"0000000000000000_0000000000000000_0000011101101110_0100111110100000"; -- 0.02902696281671524
	pesos_i(7260) := b"1111111111111111_1111111111111111_1111001010111101_0110011101100000"; -- -0.051797427237033844
	pesos_i(7261) := b"1111111111111111_1111111111111111_1110010011111000_0110101110100000"; -- -0.10558440536260605
	pesos_i(7262) := b"0000000000000000_0000000000000000_0011000000000000_1011100001000000"; -- 0.18751098215579987
	pesos_i(7263) := b"1111111111111111_1111111111111111_1100001000010111_1011000010000000"; -- -0.24182602763175964
	pesos_i(7264) := b"1111111111111111_1111111111111111_1101010011111001_1111001011000000"; -- -0.16806109249591827
	pesos_i(7265) := b"1111111111111111_1111111111111111_1101110110110001_1100111111000000"; -- -0.1340055614709854
	pesos_i(7266) := b"0000000000000000_0000000000000000_0000101010000011_1100010111100000"; -- 0.04107319563627243
	pesos_i(7267) := b"0000000000000000_0000000000000000_0001101000110001_1101010111100000"; -- 0.10232292860746384
	pesos_i(7268) := b"0000000000000000_0000000000000000_0100101100011111_0011000000000000"; -- 0.2934446334838867
	pesos_i(7269) := b"0000000000000000_0000000000000000_0000011110010001_1011111100011000"; -- 0.029567664489150047
	pesos_i(7270) := b"1111111111111111_1111111111111111_1011001010010111_1010011100000000"; -- -0.302373468875885
	pesos_i(7271) := b"0000000000000000_0000000000000000_0000110011101000_0011011001100000"; -- 0.05041828006505966
	pesos_i(7272) := b"1111111111111111_1111111111111111_1111011110000111_1100000101110000"; -- -0.03308478370308876
	pesos_i(7273) := b"0000000000000000_0000000000000000_0001001111110110_0010110010100000"; -- 0.0779750719666481
	pesos_i(7274) := b"0000000000000000_0000000000000000_0001101101011010_0001111010000000"; -- 0.10684385895729065
	pesos_i(7275) := b"1111111111111111_1111111111111111_1111000100110010_1111000011100000"; -- -0.05781645327806473
	pesos_i(7276) := b"1111111111111111_1111111111111111_1110101001011101_1000001010000000"; -- -0.08451065421104431
	pesos_i(7277) := b"1111111111111111_1111111111111111_1111100000000101_1001010001001000"; -- -0.0311648678034544
	pesos_i(7278) := b"0000000000000000_0000000000000000_0011001111100101_1010110110000000"; -- 0.20272335410118103
	pesos_i(7279) := b"1111111111111111_1111111111111111_1110110000010100_0010101001100000"; -- -0.07781729847192764
	pesos_i(7280) := b"1111111111111111_1111111111111111_1011011011011001_0101001010000000"; -- -0.28574642539024353
	pesos_i(7281) := b"0000000000000000_0000000000000000_0000010001000101_1101000010100000"; -- 0.016690291464328766
	pesos_i(7282) := b"0000000000000000_0000000000000000_0000010010010011_1000111101110000"; -- 0.01787659153342247
	pesos_i(7283) := b"0000000000000000_0000000000000000_0010110011100100_0110100101000000"; -- 0.1753602772951126
	pesos_i(7284) := b"1111111111111111_1111111111111111_1110111000010110_1101001010000000"; -- -0.06996425986289978
	pesos_i(7285) := b"0000000000000000_0000000000000000_0011000111000001_0100111101000000"; -- 0.19435591995716095
	pesos_i(7286) := b"0000000000000000_0000000000000000_0011000111101110_1001000001000000"; -- 0.19504643976688385
	pesos_i(7287) := b"1111111111111111_1111111111111111_1110111000111011_1001111100000000"; -- -0.06940275430679321
	pesos_i(7288) := b"1111111111111111_1111111111111111_1110010111001001_1100000100100000"; -- -0.10239022225141525
	pesos_i(7289) := b"1111111111111111_1111111111111111_1110101011011101_0000010100000000"; -- -0.08256500959396362
	pesos_i(7290) := b"0000000000000000_0000000000000000_0000100111001101_1001101000010000"; -- 0.03829348459839821
	pesos_i(7291) := b"0000000000000000_0000000000000000_0110010101001111_1010101000000000"; -- 0.3957468271255493
	pesos_i(7292) := b"1111111111111111_1111111111111111_1101011010011101_1100101001000000"; -- -0.16165481507778168
	pesos_i(7293) := b"0000000000000000_0000000000000000_0011001100110111_0110010000000000"; -- 0.20006394386291504
	pesos_i(7294) := b"0000000000000000_0000000000000000_0000011110111000_0110000101110000"; -- 0.030157174915075302
	pesos_i(7295) := b"0000000000000000_0000000000000000_0000110100000000_1110010010110000"; -- 0.05079488083720207
	pesos_i(7296) := b"1111111111111111_1111111111111111_0111110000010011_0111110100000000"; -- -0.5153276324272156
	pesos_i(7297) := b"0000000000000000_0000000000000000_0100000000001010_1111001100000000"; -- 0.2501670718193054
	pesos_i(7298) := b"0000000000000000_0000000000000000_0000101010111110_0000100110000000"; -- 0.041962236166000366
	pesos_i(7299) := b"1111111111111111_1111111111111111_1110100011111011_0011110110100000"; -- -0.08991637080907822
	pesos_i(7300) := b"0000000000000000_0000000000000000_0011011001000100_1011110011000000"; -- 0.21198634803295135
	pesos_i(7301) := b"1111111111111111_1111111111111111_1101001010010011_1010001110000000"; -- -0.17743471264839172
	pesos_i(7302) := b"0000000000000000_0000000000000000_0001111010010111_1111001111000000"; -- 0.1195061057806015
	pesos_i(7303) := b"0000000000000000_0000000000000000_0000000000010010_1001111010001111"; -- 0.00028410908998921514
	pesos_i(7304) := b"1111111111111111_1111111111111111_1111000101010000_1110001110100000"; -- -0.057359479367733
	pesos_i(7305) := b"1111111111111111_1111111111111111_1001100000010011_1000101100000000"; -- -0.4059517979621887
	pesos_i(7306) := b"0000000000000000_0000000000000000_0010000110010110_0010110100000000"; -- 0.1311977505683899
	pesos_i(7307) := b"0000000000000000_0000000000000000_0010110110111001_1010110000000000"; -- 0.17861437797546387
	pesos_i(7308) := b"1111111111111111_1111111111111111_1110001001111111_1011010111100000"; -- -0.11523879319429398
	pesos_i(7309) := b"0000000000000000_0000000000000000_0000001001100001_0011000111100000"; -- 0.009295575320720673
	pesos_i(7310) := b"1111111111111111_1111111111111111_1101100100000010_0100010110000000"; -- -0.1523090898990631
	pesos_i(7311) := b"0000000000000000_0000000000000000_0011111000110101_0000000001000000"; -- 0.2429962307214737
	pesos_i(7312) := b"0000000000000000_0000000000000000_0010001100000111_0010101110000000"; -- 0.13682815432548523
	pesos_i(7313) := b"0000000000000000_0000000000000000_0000111001110000_1111111001110000"; -- 0.05641165003180504
	pesos_i(7314) := b"1111111111111111_1111111111111111_1010110010100011_1001010110000000"; -- -0.3256289064884186
	pesos_i(7315) := b"1111111111111111_1111111111111111_1100110111000000_0111111100000000"; -- -0.19628149271011353
	pesos_i(7316) := b"1111111111111111_1111111111111111_1100010100010100_0111000011000000"; -- -0.23015685379505157
	pesos_i(7317) := b"0000000000000000_0000000000000000_0100000010001110_1001001000000000"; -- 0.2521754503250122
	pesos_i(7318) := b"0000000000000000_0000000000000000_0000100011101100_1111110111010000"; -- 0.034866202622652054
	pesos_i(7319) := b"0000000000000000_0000000000000000_0001111110101000_0010011011000000"; -- 0.12365953624248505
	pesos_i(7320) := b"0000000000000000_0000000000000000_0001011001010101_1101010010100000"; -- 0.08724717050790787
	pesos_i(7321) := b"0000000000000000_0000000000000000_0010100111101011_1001100000000000"; -- 0.16375112533569336
	pesos_i(7322) := b"0000000000000000_0000000000000000_0001011111001000_0000011101100000"; -- 0.09289594739675522
	pesos_i(7323) := b"0000000000000000_0000000000000000_0000010010111111_1111000000010000"; -- 0.018553737550973892
	pesos_i(7324) := b"1111111111111111_1111111111111111_1111100110000101_0100011111110000"; -- -0.02531004324555397
	pesos_i(7325) := b"1111111111111111_1111111111111111_1100010101001001_1101101111000000"; -- -0.2293417602777481
	pesos_i(7326) := b"0000000000000000_0000000000000000_0000110101000100_1000110010110000"; -- 0.05182723328471184
	pesos_i(7327) := b"0000000000000000_0000000000000000_0001111100100101_0111000000100000"; -- 0.12166500836610794
	pesos_i(7328) := b"1111111111111111_1111111111111111_1110000011010010_1100000011000000"; -- -0.12178416550159454
	pesos_i(7329) := b"0000000000000000_0000000000000000_0001001110110011_0100011100100000"; -- 0.07695431262254715
	pesos_i(7330) := b"0000000000000000_0000000000000000_0000001010001110_0100101100011000"; -- 0.009983723983168602
	pesos_i(7331) := b"1111111111111111_1111111111111111_1101101100111000_1001000000000000"; -- -0.14366817474365234
	pesos_i(7332) := b"1111111111111111_1111111111111111_1001011110101101_1000111010000000"; -- -0.407507985830307
	pesos_i(7333) := b"0000000000000000_0000000000000000_0000101110000110_1110101111110000"; -- 0.045027490705251694
	pesos_i(7334) := b"1111111111111111_1111111111111111_1101101101101001_1101101000000000"; -- -0.14291608333587646
	pesos_i(7335) := b"1111111111111111_1111111111111111_1101001001110011_1110010100000000"; -- -0.17791908979415894
	pesos_i(7336) := b"0000000000000000_0000000000000000_0110101111110110_1100110100000000"; -- 0.42173463106155396
	pesos_i(7337) := b"1111111111111111_1111111111111111_1110011101001110_0100000110100000"; -- -0.09646215289831161
	pesos_i(7338) := b"0000000000000000_0000000000000000_0000101010000000_1101011001010000"; -- 0.041028399020433426
	pesos_i(7339) := b"0000000000000000_0000000000000000_0000001111110000_1100111100111000"; -- 0.01539321057498455
	pesos_i(7340) := b"1111111111111111_1111111111111111_1111011101100000_0011111000100000"; -- -0.03368770331144333
	pesos_i(7341) := b"1111111111111111_1111111111111111_1011000011100111_1100100100000000"; -- -0.30896323919296265
	pesos_i(7342) := b"0000000000000000_0000000000000000_0000111100010011_0101000101100000"; -- 0.0588885173201561
	pesos_i(7343) := b"0000000000000000_0000000000000000_0000000000010011_0011001110011110"; -- 0.0002929935581050813
	pesos_i(7344) := b"1111111111111111_1111111111111111_1011100111010000_0110101100000000"; -- -0.27416354417800903
	pesos_i(7345) := b"0000000000000000_0000000000000000_0000111001001000_1101000100110000"; -- 0.05579860135912895
	pesos_i(7346) := b"0000000000000000_0000000000000000_0010011111111011_1010100110000000"; -- 0.15618380904197693
	pesos_i(7347) := b"0000000000000000_0000000000000000_0001001111111101_1100111010100000"; -- 0.07809153944253922
	pesos_i(7348) := b"0000000000000000_0000000000000000_0000111111111011_0101010001110000"; -- 0.06242873892188072
	pesos_i(7349) := b"1111111111111111_1111111111111111_1011110101001110_0101011110000000"; -- -0.26052334904670715
	pesos_i(7350) := b"1111111111111111_1111111111111111_1010001100110101_0010010110000000"; -- -0.3624702990055084
	pesos_i(7351) := b"0000000000000000_0000000000000000_0011100011110100_0100111111000000"; -- 0.22247789800167084
	pesos_i(7352) := b"1111111111111111_1111111111111111_1101100010100101_0110111000000000"; -- -0.1537257432937622
	pesos_i(7353) := b"0000000000000000_0000000000000000_0100100111011010_1000100000000000"; -- 0.28849077224731445
	pesos_i(7354) := b"0000000000000000_0000000000000000_0000110110010011_1000111011110000"; -- 0.05303281173110008
	pesos_i(7355) := b"1111111111111111_1111111111111111_1110011011101111_1000100100100000"; -- -0.09790747612714767
	pesos_i(7356) := b"1111111111111111_1111111111111111_1101000001010111_1111011110000000"; -- -0.1861577332019806
	pesos_i(7357) := b"1111111111111111_1111111111111111_1010110110011101_1100111000000000"; -- -0.32181084156036377
	pesos_i(7358) := b"0000000000000000_0000000000000000_0001101001000111_0111110101000000"; -- 0.10265333950519562
	pesos_i(7359) := b"1111111111111111_1111111111111111_1110110101011111_1010101001100000"; -- -0.07275900989770889
	pesos_i(7360) := b"0000000000000000_0000000000000000_0001010010001101_1001000000000000"; -- 0.08028507232666016
	pesos_i(7361) := b"0000000000000000_0000000000000000_0001110110100000_0101100010000000"; -- 0.11572793126106262
	pesos_i(7362) := b"1111111111111111_1111111111111111_1000011110111111_0101010100000000"; -- -0.4697367548942566
	pesos_i(7363) := b"1111111111111111_1111111111111111_1101011010011011_0011001010000000"; -- -0.16169437766075134
	pesos_i(7364) := b"0000000000000000_0000000000000000_0100010010101110_0011001110000000"; -- 0.26828309893608093
	pesos_i(7365) := b"1111111111111111_1111111111111111_1100101101110011_1110100010000000"; -- -0.20526263117790222
	pesos_i(7366) := b"1111111111111111_1111111111111111_1111100110011001_0010110111111000"; -- -0.02500641532242298
	pesos_i(7367) := b"0000000000000000_0000000000000000_0000001010000110_1010000000001100"; -- 0.009866717271506786
	pesos_i(7368) := b"1111111111111111_1111111111111111_1111110100000000_1011110100001000"; -- -0.011707482859492302
	pesos_i(7369) := b"0000000000000000_0000000000000000_0001000100111010_1110100111000000"; -- 0.06730519235134125
	pesos_i(7370) := b"1111111111111111_1111111111111111_1111111110101100_1010100101110101"; -- -0.0012716378550976515
	pesos_i(7371) := b"1111111111111111_1111111111111111_1110001011000100_0101101100000000"; -- -0.11419135332107544
	pesos_i(7372) := b"1111111111111111_1111111111111111_1000101101010001_1010110000000000"; -- -0.45578503608703613
	pesos_i(7373) := b"0000000000000000_0000000000000000_0011011001011110_0010110110000000"; -- 0.21237453818321228
	pesos_i(7374) := b"0000000000000000_0000000000000000_0000100001000101_1011100111010000"; -- 0.03231393173336983
	pesos_i(7375) := b"1111111111111111_1111111111111111_1101011111101011_1110011000000000"; -- -0.15655672550201416
	pesos_i(7376) := b"0000000000000000_0000000000000000_0011101100111101_0110101000000000"; -- 0.2314058542251587
	pesos_i(7377) := b"0000000000000000_0000000000000000_0011100111111000_0111111101000000"; -- 0.22644801437854767
	pesos_i(7378) := b"1111111111111111_1111111111111111_1011110010110101_0101011100000000"; -- -0.26285797357559204
	pesos_i(7379) := b"1111111111111111_1111111111111111_1100000100011001_1000001001000000"; -- -0.2457045167684555
	pesos_i(7380) := b"1111111111111111_1111111111111111_1111101001110010_1101110100011000"; -- -0.02168481983244419
	pesos_i(7381) := b"0000000000000000_0000000000000000_0101010111100001_1101100100000000"; -- 0.33547741174697876
	pesos_i(7382) := b"0000000000000000_0000000000000000_0011110110110110_0110111110000000"; -- 0.24106499552726746
	pesos_i(7383) := b"0000000000000000_0000000000000000_0010000110110011_1100011111000000"; -- 0.13164947926998138
	pesos_i(7384) := b"0000000000000000_0000000000000000_0111110100110111_0000100010000000"; -- 0.4891209900379181
	pesos_i(7385) := b"0000000000000000_0000000000000000_0001001110110011_0001101101100000"; -- 0.07695170491933823
	pesos_i(7386) := b"1111111111111111_1111111111111111_1111101111001010_1111101101011000"; -- -0.016433993354439735
	pesos_i(7387) := b"0000000000000000_0000000000000000_0001010110001101_0111001011000000"; -- 0.08418957889080048
	pesos_i(7388) := b"0000000000000000_0000000000000000_0001110011011110_1001010011000000"; -- 0.11277131736278534
	pesos_i(7389) := b"1111111111111111_1111111111111111_1110100110001101_1110110011000000"; -- -0.08767814934253693
	pesos_i(7390) := b"0000000000000000_0000000000000000_0010111111010010_0100100011000000"; -- 0.1868024319410324
	pesos_i(7391) := b"1111111111111111_1111111111111111_1110010011110101_0011001100000000"; -- -0.10563355684280396
	pesos_i(7392) := b"1111111111111111_1111111111111111_1100000001101011_1001010100000000"; -- -0.24835842847824097
	pesos_i(7393) := b"0000000000000000_0000000000000000_0000000100101100_0110110011100000"; -- 0.004584126174449921
	pesos_i(7394) := b"0000000000000000_0000000000000000_0011101110011110_0000010011000000"; -- 0.23287992179393768
	pesos_i(7395) := b"0000000000000000_0000000000000000_1000100111000101_0111001000000000"; -- 0.5381690263748169
	pesos_i(7396) := b"0000000000000000_0000000000000000_0011000011111011_0110001001000000"; -- 0.19133581221103668
	pesos_i(7397) := b"1111111111111111_1111111111111111_1101000101110100_1110111100000000"; -- -0.18180948495864868
	pesos_i(7398) := b"1111111111111111_1111111111111111_1010100100111100_1011110100000000"; -- -0.33891695737838745
	pesos_i(7399) := b"1111111111111111_1111111111111111_1111001000010011_0000101110100000"; -- -0.054396890103816986
	pesos_i(7400) := b"0000000000000000_0000000000000000_0011010110001100_1011100001000000"; -- 0.20917846262454987
	pesos_i(7401) := b"0000000000000000_0000000000000000_0001111111001000_1011011100000000"; -- 0.1241564154624939
	pesos_i(7402) := b"0000000000000000_0000000000000000_0110000001111100_1100110010000000"; -- 0.37690427899360657
	pesos_i(7403) := b"1111111111111111_1111111111111111_1010000101001000_1011001010000000"; -- -0.3699844777584076
	pesos_i(7404) := b"0000000000000000_0000000000000000_0000001010011100_0111111101101000"; -- 0.010200465098023415
	pesos_i(7405) := b"0000000000000000_0000000000000000_0110111011111101_1111111010000000"; -- 0.43356314301490784
	pesos_i(7406) := b"1111111111111111_1111111111111111_1101001001111011_0010000110000000"; -- -0.17780867218971252
	pesos_i(7407) := b"1111111111111111_1111111111111111_1101000101110110_1000100100000000"; -- -0.18178504705429077
	pesos_i(7408) := b"1111111111111111_1111111111111111_1001001000111101_0011100010000000"; -- -0.4287533462047577
	pesos_i(7409) := b"1111111111111111_1111111111111111_1111100001000100_0011011001100000"; -- -0.030209161341190338
	pesos_i(7410) := b"0000000000000000_0000000000000000_0001111100010011_0110011111100000"; -- 0.12138985842466354
	pesos_i(7411) := b"0000000000000000_0000000000000000_0010101010001011_1000101100000000"; -- 0.16619175672531128
	pesos_i(7412) := b"1111111111111111_1111111111111111_1100001110000011_0011101110000000"; -- -0.23627880215644836
	pesos_i(7413) := b"1111111111111111_1111111111111111_1011110111110001_1100110010000000"; -- -0.25802919268608093
	pesos_i(7414) := b"0000000000000000_0000000000000000_0010110110110011_0000111111000000"; -- 0.1785135120153427
	pesos_i(7415) := b"0000000000000000_0000000000000000_0001111010001011_0000100011000000"; -- 0.11930899322032928
	pesos_i(7416) := b"1111111111111111_1111111111111111_1110010010011111_0100011001000000"; -- -0.10694466531276703
	pesos_i(7417) := b"0000000000000000_0000000000000000_0011000100010101_0110101100000000"; -- 0.19173306226730347
	pesos_i(7418) := b"1111111111111111_1111111111111111_1111100001011011_0101110110110000"; -- -0.029855865985155106
	pesos_i(7419) := b"0000000000000000_0000000000000000_0011100111011110_0101110110000000"; -- 0.2260492742061615
	pesos_i(7420) := b"0000000000000000_0000000000000000_0010110101101010_0000000110000000"; -- 0.17739877104759216
	pesos_i(7421) := b"1111111111111111_1111111111111111_1111001110101101_0111000100010000"; -- -0.04813474044203758
	pesos_i(7422) := b"0000000000000000_0000000000000000_0001111000011110_1101111010100000"; -- 0.11765853315591812
	pesos_i(7423) := b"0000000000000000_0000000000000000_0011111010111000_0010111100000000"; -- 0.24499791860580444
	pesos_i(7424) := b"1111111111111111_1111111111111111_0101100101001101_0110010000000000"; -- -0.65116286277771
	pesos_i(7425) := b"0000000000000000_0000000000000000_0101110001001110_0011100000000000"; -- 0.3605685234069824
	pesos_i(7426) := b"0000000000000000_0000000000000000_0010010111001111_0001010001000000"; -- 0.1476910263299942
	pesos_i(7427) := b"1111111111111111_1111111111111111_1111110000100111_1111011001110000"; -- -0.015015218406915665
	pesos_i(7428) := b"0000000000000000_0000000000000000_0100001101001110_1100000000000000"; -- 0.2629203796386719
	pesos_i(7429) := b"1111111111111111_1111111111111111_1100011101111001_0010110010000000"; -- -0.220807284116745
	pesos_i(7430) := b"0000000000000000_0000000000000000_0010111111101001_1101111100000000"; -- 0.1871623396873474
	pesos_i(7431) := b"0000000000000000_0000000000000000_0011001001011011_0000110001000000"; -- 0.196701779961586
	pesos_i(7432) := b"1111111111111111_1111111111111111_1110010101111110_1000000101000000"; -- -0.10353843867778778
	pesos_i(7433) := b"1111111111111111_1111111111111111_1011001101000101_1110110100000000"; -- -0.29971426725387573
	pesos_i(7434) := b"0000000000000000_0000000000000000_0110010100110101_1110011100000000"; -- 0.3953537344932556
	pesos_i(7435) := b"0000000000000000_0000000000000000_0001010010001110_1011110011000000"; -- 0.08030299842357635
	pesos_i(7436) := b"1111111111111111_1111111111111111_1110100010101000_1100001100100000"; -- -0.0911748930811882
	pesos_i(7437) := b"1111111111111111_1111111111111111_0111100010101010_0010011000000000"; -- -0.5286537408828735
	pesos_i(7438) := b"1111111111111111_1111111111111111_0010101011011010_1001001000000000"; -- -0.8326023817062378
	pesos_i(7439) := b"0000000000000000_0000000000000000_0100101011110010_1010101010000000"; -- 0.2927652895450592
	pesos_i(7440) := b"1111111111111111_1111111111111111_1111001101110001_0011100100110000"; -- -0.04905359819531441
	pesos_i(7441) := b"1111111111111111_1111111111111111_1111000100101001_0101000001010000"; -- -0.057963352650403976
	pesos_i(7442) := b"1111111111111111_1111111111111111_1001011111100001_1001110010000000"; -- -0.40671369433403015
	pesos_i(7443) := b"1111111111111111_1111111111111111_0111101011010100_0101101100000000"; -- -0.5201972126960754
	pesos_i(7444) := b"1111111111111111_1111111111111111_1111100100010010_1111111110001000"; -- -0.02705386094748974
	pesos_i(7445) := b"1111111111111111_1111111111111111_1111111110100001_1101110111010110"; -- -0.0014363625086843967
	pesos_i(7446) := b"0000000000000000_0000000000000000_0100110101001000_1001000010000000"; -- 0.30188849568367004
	pesos_i(7447) := b"0000000000000000_0000000000000000_0001111100010111_0100011010100000"; -- 0.12144891172647476
	pesos_i(7448) := b"0000000000000000_0000000000000000_0000010101110000_0101000101011000"; -- 0.021245082840323448
	pesos_i(7449) := b"0000000000000000_0000000000000000_0100011011011010_0101001110000000"; -- 0.27676889300346375
	pesos_i(7450) := b"1111111111111111_1111111111111111_1111010111101010_1000001100010000"; -- -0.039390381425619125
	pesos_i(7451) := b"0000000000000000_0000000000000000_0001010101011101_0011001111100000"; -- 0.08345340937376022
	pesos_i(7452) := b"1111111111111111_1111111111111111_1110100100011101_1000000110000000"; -- -0.08939352631568909
	pesos_i(7453) := b"1111111111111111_1111111111111111_1110111011100111_0001101011000000"; -- -0.06678612530231476
	pesos_i(7454) := b"0000000000000000_0000000000000000_0001010111011011_0110101111000000"; -- 0.08537934720516205
	pesos_i(7455) := b"0000000000000000_0000000000000000_0000001110101000_0111100101010000"; -- 0.014289457350969315
	pesos_i(7456) := b"1111111111111111_1111111111111111_1111011100010000_1111010010100000"; -- -0.03489752858877182
	pesos_i(7457) := b"1111111111111111_1111111111111111_1001101001011101_0000110100000000"; -- -0.3970176577568054
	pesos_i(7458) := b"0000000000000000_0000000000000000_0000101001111010_0011000001000000"; -- 0.04092694818973541
	pesos_i(7459) := b"0000000000000000_0000000000000000_0010101010101000_0111010110000000"; -- 0.1666329801082611
	pesos_i(7460) := b"1111111111111111_1111111111111111_1001001100001000_1111001110000000"; -- -0.4256446659564972
	pesos_i(7461) := b"1111111111111111_1111111111111111_1111101101111000_1100100010111000"; -- -0.01768823154270649
	pesos_i(7462) := b"0000000000000000_0000000000000000_0001010101101010_0011100100100000"; -- 0.0836520865559578
	pesos_i(7463) := b"1111111111111111_1111111111111111_1101101010100110_0110110010000000"; -- -0.14589807391166687
	pesos_i(7464) := b"0000000000000000_0000000000000000_1001010101000100_0101011000000000"; -- 0.5830739736557007
	pesos_i(7465) := b"1111111111111111_1111111111111111_1110000010101100_1001010110100000"; -- -0.12236656993627548
	pesos_i(7466) := b"1111111111111111_1111111111111111_1100010101001111_0110101110000000"; -- -0.22925689816474915
	pesos_i(7467) := b"0000000000000000_0000000000000000_0011001001111010_1000100110000000"; -- 0.19718226790428162
	pesos_i(7468) := b"0000000000000000_0000000000000000_0000101001101111_0111101100100000"; -- 0.04076356440782547
	pesos_i(7469) := b"1111111111111111_1111111111111111_1101101111111011_1100011000000000"; -- -0.14068949222564697
	pesos_i(7470) := b"0000000000000000_0000000000000000_0110110111101011_1100011010000000"; -- 0.4293788969516754
	pesos_i(7471) := b"0000000000000000_0000000000000000_0001101001011000_1001011010100000"; -- 0.1029142513871193
	pesos_i(7472) := b"1111111111111111_1111111111111111_1010100000011111_1011001110000000"; -- -0.3432662785053253
	pesos_i(7473) := b"1111111111111111_1111111111111111_1010111010101011_1110011010000000"; -- -0.3176895081996918
	pesos_i(7474) := b"0000000000000000_0000000000000000_0101101100110001_0011001100000000"; -- 0.35621947050094604
	pesos_i(7475) := b"1111111111111111_1111111111111111_1100011101111000_0110011110000000"; -- -0.22081902623176575
	pesos_i(7476) := b"0000000000000000_0000000000000000_0100001111001001_1100011110000000"; -- 0.2647976577281952
	pesos_i(7477) := b"1111111111111111_1111111111111111_1110111100110101_0001001010000000"; -- -0.06559643149375916
	pesos_i(7478) := b"1111111111111111_1111111111111111_1101011000111101_1011110100000000"; -- -0.16312044858932495
	pesos_i(7479) := b"0000000000000000_0000000000000000_1000110110000111_0101000000000000"; -- 0.5528459548950195
	pesos_i(7480) := b"1111111111111111_1111111111111111_1101100011111111_0100001101000000"; -- -0.15235500037670135
	pesos_i(7481) := b"1111111111111111_1111111111111111_1100101111001100_0101011000000000"; -- -0.20391333103179932
	pesos_i(7482) := b"0000000000000000_0000000000000000_0100100000000011_1100001000000000"; -- 0.2813073396682739
	pesos_i(7483) := b"0000000000000000_0000000000000000_0001000111100110_0001110011100000"; -- 0.06991749256849289
	pesos_i(7484) := b"1111111111111111_1111111111111111_1110111000001011_0110111111100000"; -- -0.07013798505067825
	pesos_i(7485) := b"1111111111111111_1111111111111111_1000111101000100_0110110000000000"; -- -0.44036221504211426
	pesos_i(7486) := b"0000000000000000_0000000000000000_0100000100001001_1101110110000000"; -- 0.25405678153038025
	pesos_i(7487) := b"1111111111111111_1111111111111111_1100101001001000_0001011000000000"; -- -0.20983755588531494
	pesos_i(7488) := b"0000000000000000_0000000000000000_0010010100001011_1001011110000000"; -- 0.14470812678337097
	pesos_i(7489) := b"0000000000000000_0000000000000000_0100000010101100_1011001000000000"; -- 0.25263512134552
	pesos_i(7490) := b"1111111111111111_1111111111111111_1100000100110110_0010101101000000"; -- -0.24526719748973846
	pesos_i(7491) := b"1111111111111111_1111111111111111_1110011100001011_1010011111100000"; -- -0.09747839719057083
	pesos_i(7492) := b"0000000000000000_0000000000000000_0100000110100101_1000001000000000"; -- 0.2564316987991333
	pesos_i(7493) := b"1111111111111111_1111111111111111_1011001000111000_1010011000000000"; -- -0.3038231134414673
	pesos_i(7494) := b"0000000000000000_0000000000000000_0010000001100111_1100101110000000"; -- 0.1265837848186493
	pesos_i(7495) := b"0000000000000000_0000000000000000_0011011001011001_0111111111000000"; -- 0.21230314671993256
	pesos_i(7496) := b"1111111111111111_1111111111111111_0111010111111001_1000000100000000"; -- -0.5391616225242615
	pesos_i(7497) := b"0000000000000000_0000000000000000_0000001010100110_0010011111100100"; -- 0.010347836650907993
	pesos_i(7498) := b"0000000000000000_0000000000000000_0011011011010000_0100111100000000"; -- 0.21411603689193726
	pesos_i(7499) := b"1111111111111111_1111111111111111_1000000101101001_0001101000000000"; -- -0.49449002742767334
	pesos_i(7500) := b"1111111111111111_1111111111111111_1001100000101111_0010100000000000"; -- -0.4055304527282715
	pesos_i(7501) := b"0000000000000000_0000000000000000_0111110000101010_1011011010000000"; -- 0.4850267469882965
	pesos_i(7502) := b"0000000000000000_0000000000000000_0001010101011101_0101010010100000"; -- 0.08345536142587662
	pesos_i(7503) := b"1111111111111111_1111111111111111_1110011000010111_1011111110100000"; -- -0.10120012611150742
	pesos_i(7504) := b"0000000000000000_0000000000000000_0100000111110100_0011011000000000"; -- 0.25763261318206787
	pesos_i(7505) := b"0000000000000000_0000000000000000_0110011011010101_1101110110000000"; -- 0.40170082449913025
	pesos_i(7506) := b"1111111111111111_1111111111111111_1000010010001001_0001110000000000"; -- -0.4822828769683838
	pesos_i(7507) := b"1111111111111111_1111111111111111_1011011000001100_1101101010000000"; -- -0.2888663709163666
	pesos_i(7508) := b"0000000000000000_0000000000000000_0010000110011011_1011000011000000"; -- 0.13128189742565155
	pesos_i(7509) := b"0000000000000000_0000000000000000_1000111011001011_1100011100000000"; -- 0.5577968955039978
	pesos_i(7510) := b"0000000000000000_0000000000000000_0101110000011011_0001010100000000"; -- 0.3597882390022278
	pesos_i(7511) := b"0000000000000000_0000000000000000_0010000001010111_0100110010000000"; -- 0.12633207440376282
	pesos_i(7512) := b"0000000000000000_0000000000000000_1001000001010001_0110010000000000"; -- 0.56374192237854
	pesos_i(7513) := b"0000000000000000_0000000000000000_0100000111101110_0010000110000000"; -- 0.257539838552475
	pesos_i(7514) := b"0000000000000000_0000000000000000_0011010111100111_0110101100000000"; -- 0.21056240797042847
	pesos_i(7515) := b"1111111111111111_1111111111111111_1111011000101110_1000001100010000"; -- -0.038352783769369125
	pesos_i(7516) := b"0000000000000000_0000000000000000_0010000011001111_1000001111000000"; -- 0.12816642224788666
	pesos_i(7517) := b"0000000000000000_0000000000000000_0000100111101110_1111000110000000"; -- 0.03880223631858826
	pesos_i(7518) := b"0000000000000000_0000000000000000_0111101100110100_1100101100000000"; -- 0.4812743067741394
	pesos_i(7519) := b"0000000000000000_0000000000000000_0000001110110000_0100101101011100"; -- 0.01440878864377737
	pesos_i(7520) := b"1111111111111111_1111111111111111_1011010110111010_0011111010000000"; -- -0.29012688994407654
	pesos_i(7521) := b"0000000000000000_0000000000000000_0000011101010001_1110010010000000"; -- 0.028593331575393677
	pesos_i(7522) := b"0000000000000000_0000000000000000_0110000101001100_1011010000000000"; -- 0.38007664680480957
	pesos_i(7523) := b"0000000000000000_0000000000000000_1011000010101110_1101100100000000"; -- 0.6901679635047913
	pesos_i(7524) := b"0000000000000000_0000000000000000_0110110100001100_0000101010000000"; -- 0.42596498131752014
	pesos_i(7525) := b"1111111111111111_1111111111111111_1100101011101111_1111011111000000"; -- -0.2072758823633194
	pesos_i(7526) := b"1111111111111111_1111111111111111_1011110101000011_0001111010000000"; -- -0.26069459319114685
	pesos_i(7527) := b"1111111111111111_1111111111111111_1010101100100001_0101101100000000"; -- -0.33152228593826294
	pesos_i(7528) := b"0000000000000000_0000000000000000_0011001101000010_0110100111000000"; -- 0.20023213326931
	pesos_i(7529) := b"1111111111111111_1111111111111111_1111010110000001_1110110000000000"; -- -0.04098629951477051
	pesos_i(7530) := b"0000000000000000_0000000000000000_1000011110100100_0010011100000000"; -- 0.5298485159873962
	pesos_i(7531) := b"1111111111111111_1111111111111111_0101000101100101_0011010000000000"; -- -0.6820495128631592
	pesos_i(7532) := b"1111111111111111_1111111111111111_1110000011000110_1101011000100000"; -- -0.12196599692106247
	pesos_i(7533) := b"0000000000000000_0000000000000000_0001010111001110_0110010000000000"; -- 0.08518052101135254
	pesos_i(7534) := b"1111111111111111_1111111111111111_1101101110101001_1000100100000000"; -- -0.14194434881210327
	pesos_i(7535) := b"1111111111111111_1111111111111111_1100010101100100_0011010110000000"; -- -0.22893968224525452
	pesos_i(7536) := b"1111111111111111_1111111111111111_0110100100000010_1010001000000000"; -- -0.5898035764694214
	pesos_i(7537) := b"1111111111111111_1111111111111111_1011001111000001_0011001110000000"; -- -0.29783323407173157
	pesos_i(7538) := b"0000000000000000_0000000000000000_0000011111010011_1110010000001000"; -- 0.03057694621384144
	pesos_i(7539) := b"0000000000000000_0000000000000000_0101100111000000_1010110110000000"; -- 0.35059627890586853
	pesos_i(7540) := b"1111111111111111_1111111111111111_1100011110000111_1000000111000000"; -- -0.2205885797739029
	pesos_i(7541) := b"1111111111111111_1111111111111111_1111100100111111_1000101110110000"; -- -0.026374120265245438
	pesos_i(7542) := b"1111111111111111_1111111111111111_1111000000001000_1100100111000000"; -- -0.062365904450416565
	pesos_i(7543) := b"0000000000000000_0000000000000000_0001010000100001_0110000011000000"; -- 0.07863430678844452
	pesos_i(7544) := b"1111111111111111_1111111111111111_1001000101000011_0011001010000000"; -- -0.43256840109825134
	pesos_i(7545) := b"0000000000000000_0000000000000000_0010000100101010_1101110000000000"; -- 0.12956023216247559
	pesos_i(7546) := b"1111111111111111_1111111111111111_1100011000010110_0110000110000000"; -- -0.2262209951877594
	pesos_i(7547) := b"0000000000000000_0000000000000000_1001110000100011_0011100000000000"; -- 0.6099123954772949
	pesos_i(7548) := b"0000000000000000_0000000000000000_0011110000100001_0010100010000000"; -- 0.2348809540271759
	pesos_i(7549) := b"0000000000000000_0000000000000000_0011001011101110_0010000100000000"; -- 0.1989460587501526
	pesos_i(7550) := b"1111111111111111_1111111111111111_1111011010100110_1000101011110000"; -- -0.03652125969529152
	pesos_i(7551) := b"0000000000000000_0000000000000000_0100101000000011_0000110000000000"; -- 0.2891089916229248
	pesos_i(7552) := b"1111111111111111_1111111111111111_1111010000110011_0011011000000000"; -- -0.04609358310699463
	pesos_i(7553) := b"0000000000000000_0000000000000000_1010111101001011_0010110000000000"; -- 0.6847407817840576
	pesos_i(7554) := b"0000000000000000_0000000000000000_0000000000101110_0001101100111100"; -- 0.0007035275339148939
	pesos_i(7555) := b"1111111111111111_1111111111111111_1111001100101000_1000110001010000"; -- -0.05016253516077995
	pesos_i(7556) := b"0000000000000000_0000000000000000_0010100010011011_1110111011000000"; -- 0.15862934291362762
	pesos_i(7557) := b"0000000000000000_0000000000000000_0000001100000011_0010101111011000"; -- 0.011767139658331871
	pesos_i(7558) := b"0000000000000000_0000000000000000_0000110010000011_0101100101000000"; -- 0.048879221081733704
	pesos_i(7559) := b"1111111111111111_1111111111111111_1011011101011011_0000011000000000"; -- -0.28376734256744385
	pesos_i(7560) := b"0000000000000000_0000000000000000_0010101100010101_1111100000000000"; -- 0.1683039665222168
	pesos_i(7561) := b"1111111111111111_1111111111111111_1110001000100111_0001011001000000"; -- -0.11659108102321625
	pesos_i(7562) := b"0000000000000000_0000000000000000_1011010111001001_0011001000000000"; -- 0.7101012468338013
	pesos_i(7563) := b"0000000000000000_0000000000000000_0101001101100011_1100000000000000"; -- 0.3257408142089844
	pesos_i(7564) := b"1111111111111111_1111111111111111_1001000100011011_0000101100000000"; -- -0.43318110704421997
	pesos_i(7565) := b"1111111111111111_1111111111111111_0100100110101110_1011101000000000"; -- -0.7121776342391968
	pesos_i(7566) := b"1111111111111111_1111111111111110_1110000111011010_1000111000000000"; -- -1.117758870124817
	pesos_i(7567) := b"0000000000000000_0000000000000000_0110010111010101_0001101110000000"; -- 0.3977830111980438
	pesos_i(7568) := b"0000000000000000_0000000000000000_0001100100001001_1001011010000000"; -- 0.0978025496006012
	pesos_i(7569) := b"0000000000000000_0000000000000000_0000110010000111_1010001010110000"; -- 0.048944633454084396
	pesos_i(7570) := b"1111111111111111_1111111111111111_1110001001111001_0101110011000000"; -- -0.11533565819263458
	pesos_i(7571) := b"1111111111111111_1111111111111111_1010010010011001_0100001010000000"; -- -0.35703644156455994
	pesos_i(7572) := b"0000000000000000_0000000000000000_0001000011011011_0101001110000000"; -- 0.06584665179252625
	pesos_i(7573) := b"1111111111111111_1111111111111111_1110000101010111_0001101010100000"; -- -0.11976464837789536
	pesos_i(7574) := b"0000000000000000_0000000000000000_0101111110101101_0110000010000000"; -- 0.3737392723560333
	pesos_i(7575) := b"0000000000000000_0000000000000000_0011010011001011_1001001000000000"; -- 0.2062312364578247
	pesos_i(7576) := b"1111111111111111_1111111111111111_1101111010001001_0111001000000000"; -- -0.1307152509689331
	pesos_i(7577) := b"0000000000000000_0000000000000000_0101100011100111_1111101100000000"; -- 0.3472897410392761
	pesos_i(7578) := b"0000000000000000_0000000000000000_0110011100010011_1011100110000000"; -- 0.40264472365379333
	pesos_i(7579) := b"0000000000000000_0000000000000000_0100001100100101_1110110100000000"; -- 0.26229745149612427
	pesos_i(7580) := b"1111111111111111_1111111111111111_1100111001100001_0011000111000000"; -- -0.19382943212985992
	pesos_i(7581) := b"1111111111111111_1111111111111111_1110110110011001_0100110110000000"; -- -0.07187953591346741
	pesos_i(7582) := b"0000000000000000_0000000000000000_1001110010111010_1111110000000000"; -- 0.6122281551361084
	pesos_i(7583) := b"0000000000000000_0000000000000000_0010101110001011_1110110000000000"; -- 0.1701037883758545
	pesos_i(7584) := b"1111111111111111_1111111111111111_1001110101110111_0101111000000000"; -- -0.3848973512649536
	pesos_i(7585) := b"1111111111111111_1111111111111111_0110110111101110_0000100100000000"; -- -0.570586621761322
	pesos_i(7586) := b"0000000000000000_0000000000000000_0100111001101110_1001000110000000"; -- 0.3063746392726898
	pesos_i(7587) := b"0000000000000000_0000000000000000_0010010101010000_0111010011000000"; -- 0.14575891196727753
	pesos_i(7588) := b"1111111111111111_1111111111111111_0110011001001101_1101001000000000"; -- -0.6003750562667847
	pesos_i(7589) := b"0000000000000000_0000000000000000_0010001110111001_0100011100000000"; -- 0.13954585790634155
	pesos_i(7590) := b"1111111111111111_1111111111111111_1111101110001011_1100010100010000"; -- -0.01739853248000145
	pesos_i(7591) := b"0000000000000000_0000000000000000_0010011011100010_0101100000000000"; -- 0.15189123153686523
	pesos_i(7592) := b"0000000000000000_0000000000000000_0101010100100011_1010110000000000"; -- 0.33257555961608887
	pesos_i(7593) := b"1111111111111111_1111111111111111_1111000100010110_0100000100010000"; -- -0.0582541786134243
	pesos_i(7594) := b"1111111111111111_1111111111111111_1111000001111000_1101000101000000"; -- -0.06065647304058075
	pesos_i(7595) := b"1111111111111111_1111111111111111_1110001010000011_1001000111000000"; -- -0.11517991125583649
	pesos_i(7596) := b"0000000000000000_0000000000000000_0010001000010000_0011111111000000"; -- 0.13306044042110443
	pesos_i(7597) := b"0000000000000000_0000000000000000_0010110001011010_0000100001000000"; -- 0.1732487827539444
	pesos_i(7598) := b"0000000000000000_0000000000000000_0110101010000010_0001110010000000"; -- 0.4160478413105011
	pesos_i(7599) := b"0000000000000000_0000000000000000_0011110110110111_0010100011000000"; -- 0.2410760372877121
	pesos_i(7600) := b"0000000000000000_0000000000000000_0001001101100100_0111001111000000"; -- 0.07575152814388275
	pesos_i(7601) := b"1111111111111111_1111111111111111_1011110110000110_1010001000000000"; -- -0.2596644163131714
	pesos_i(7602) := b"0000000000000000_0000000000000000_0000111101010001_0001110010110000"; -- 0.059831421822309494
	pesos_i(7603) := b"1111111111111111_1111111111111111_1111110000001000_1001111000010000"; -- -0.01549350842833519
	pesos_i(7604) := b"0000000000000000_0000000000000000_0010100010111001_1100101011000000"; -- 0.1590849608182907
	pesos_i(7605) := b"0000000000000000_0000000000000000_0001000100001010_1101011011000000"; -- 0.06657163798809052
	pesos_i(7606) := b"0000000000000000_0000000000000000_0010011110110010_0100000101000000"; -- 0.1550637036561966
	pesos_i(7607) := b"0000000000000000_0000000000000000_1101101101001101_1000000100000000"; -- 0.8566513657569885
	pesos_i(7608) := b"0000000000000000_0000000000000000_0000100000001101_1110110110000000"; -- 0.031462520360946655
	pesos_i(7609) := b"0000000000000000_0000000000000000_0110111101110010_1001011010000000"; -- 0.4353422224521637
	pesos_i(7610) := b"0000000000000000_0000000000000000_0000110011001011_1110001000000000"; -- 0.04998600482940674
	pesos_i(7611) := b"0000000000000000_0000000000000000_0110101111010110_0101010100000000"; -- 0.4212391972541809
	pesos_i(7612) := b"0000000000000000_0000000000000000_0100110011101011_0000011000000000"; -- 0.30046117305755615
	pesos_i(7613) := b"1111111111111111_1111111111111111_1101101010110001_0111101101000000"; -- -0.14572934806346893
	pesos_i(7614) := b"0000000000000000_0000000000000000_0101101111100110_1111000110000000"; -- 0.35899266600608826
	pesos_i(7615) := b"1111111111111111_1111111111111111_0011100111011000_1010010100000000"; -- -0.7740380167961121
	pesos_i(7616) := b"1111111111111111_1111111111111111_1101111011001000_1000101011000000"; -- -0.12975247204303741
	pesos_i(7617) := b"1111111111111111_1111111111111111_1011010110000010_1010110000000000"; -- -0.29097485542297363
	pesos_i(7618) := b"0000000000000000_0000000000000000_0100001000111110_1000010000000000"; -- 0.25876641273498535
	pesos_i(7619) := b"0000000000000000_0000000000000000_0010000101111001_1110111110000000"; -- 0.1307668387889862
	pesos_i(7620) := b"0000000000000000_0000000000000000_0101001011010100_1010000000000000"; -- 0.32355690002441406
	pesos_i(7621) := b"1111111111111111_1111111111111111_1111010111001001_0101001000010000"; -- -0.03989684209227562
	pesos_i(7622) := b"0000000000000000_0000000000000000_0111100010101010_0010100010000000"; -- 0.4713464081287384
	pesos_i(7623) := b"0000000000000000_0000000000000000_0011011010101001_1110100101000000"; -- 0.21353013813495636
	pesos_i(7624) := b"1111111111111111_1111111111111111_0110000011010001_1100010100000000"; -- -0.6217991709709167
	pesos_i(7625) := b"0000000000000000_0000000000000000_0100101000110100_0011000110000000"; -- 0.2898589074611664
	pesos_i(7626) := b"1111111111111111_1111111111111111_1111011001010101_0111001110010000"; -- -0.037758614867925644
	pesos_i(7627) := b"1111111111111111_1111111111111111_0011111100011010_0100101100000000"; -- -0.7535050511360168
	pesos_i(7628) := b"1111111111111111_1111111111111111_1110010000011001_0001010110100000"; -- -0.10899224132299423
	pesos_i(7629) := b"0000000000000000_0000000000000000_1001011001110111_1111001000000000"; -- 0.5877677202224731
	pesos_i(7630) := b"1111111111111111_1111111111111111_1000111101011110_1000100110000000"; -- -0.4399637281894684
	pesos_i(7631) := b"1111111111111111_1111111111111111_1110000110100010_1011010001000000"; -- -0.11861108243465424
	pesos_i(7632) := b"0000000000000000_0000000000000000_0001010010110000_1000001000000000"; -- 0.0808182954788208
	pesos_i(7633) := b"0000000000000000_0000000000000000_0000101100111010_0010011010100000"; -- 0.04385606199502945
	pesos_i(7634) := b"1111111111111111_1111111111111111_0111110001111000_0010011000000000"; -- -0.5137916803359985
	pesos_i(7635) := b"1111111111111111_1111111111111111_0111111111111011_0001000100000000"; -- -0.5000752806663513
	pesos_i(7636) := b"0000000000000000_0000000000000000_0101010101110011_0101001000000000"; -- 0.3337908983230591
	pesos_i(7637) := b"0000000000000000_0000000000000000_0101111111011000_1001001010000000"; -- 0.3743983805179596
	pesos_i(7638) := b"1111111111111111_1111111111111111_1101001111101101_0110011000000000"; -- -0.1721588373184204
	pesos_i(7639) := b"0000000000000000_0000000000000000_0010111000111110_1000111100000000"; -- 0.18064206838607788
	pesos_i(7640) := b"0000000000000000_0000000000000000_1001111010101100_0010001100000000"; -- 0.6198140978813171
	pesos_i(7641) := b"1111111111111111_1111111111111111_1100111010010100_0011011001000000"; -- -0.19305096566677094
	pesos_i(7642) := b"1111111111111111_1111111111111111_1111100000101111_1110000010010000"; -- -0.030519451946020126
	pesos_i(7643) := b"0000000000000000_0000000000000000_0000001001001000_0111101111001100"; -- 0.008918511681258678
	pesos_i(7644) := b"1111111111111111_1111111111111111_1110100111100011_0100111110100000"; -- -0.08637525886297226
	pesos_i(7645) := b"0000000000000000_0000000000000000_0000001101101011_1001001001011100"; -- 0.013360164128243923
	pesos_i(7646) := b"0000000000000000_0000000000000000_1010011101000000_1101101100000000"; -- 0.6533333659172058
	pesos_i(7647) := b"1111111111111111_1111111111111111_1011100101001110_0010101010000000"; -- -0.27615103125572205
	pesos_i(7648) := b"0000000000000000_0000000000000000_0101100110011000_0011110010000000"; -- 0.3499791920185089
	pesos_i(7649) := b"1111111111111111_1111111111111111_1110011111100000_0010111110000000"; -- -0.09423545002937317
	pesos_i(7650) := b"0000000000000000_0000000000000000_0110110100111110_0011100110000000"; -- 0.4267307221889496
	pesos_i(7651) := b"0000000000000000_0000000000000000_0111101001101100_1110111010000000"; -- 0.47822466492652893
	pesos_i(7652) := b"0000000000000000_0000000000000000_1001101111000010_1100011100000000"; -- 0.6084408164024353
	pesos_i(7653) := b"1111111111111111_1111111111111111_1011011111110110_0100000110000000"; -- -0.2813986837863922
	pesos_i(7654) := b"1111111111111111_1111111111111111_1100010111010101_1100111110000000"; -- -0.2272062599658966
	pesos_i(7655) := b"1111111111111111_1111111111111111_1110010001111011_0111100001100000"; -- -0.10749099403619766
	pesos_i(7656) := b"0000000000000000_0000000000000000_0000011001011011_1011110010010000"; -- 0.02483728900551796
	pesos_i(7657) := b"1111111111111111_1111111111111111_1011101000001001_0000000010000000"; -- -0.2733001410961151
	pesos_i(7658) := b"0000000000000000_0000000000000000_1101001100100011_0100011000000000"; -- 0.8247569799423218
	pesos_i(7659) := b"1111111111111111_1111111111111111_0011111101010101_1110001100000000"; -- -0.7525957226753235
	pesos_i(7660) := b"1111111111111111_1111111111111111_1011010101111100_0001010100000000"; -- -0.2910754084587097
	pesos_i(7661) := b"0000000000000000_0000000000000000_0001110010010000_0011110101000000"; -- 0.11157591640949249
	pesos_i(7662) := b"0000000000000000_0000000000000000_0001000000111100_0111111000000000"; -- 0.0634230375289917
	pesos_i(7663) := b"0000000000000000_0000000000000000_0010101010110010_0011100110000000"; -- 0.16678199172019958
	pesos_i(7664) := b"1111111111111111_1111111111111111_0110001001001110_1100011000000000"; -- -0.6159855127334595
	pesos_i(7665) := b"1111111111111111_1111111111111111_1000100000010011_1001011010000000"; -- -0.4684511125087738
	pesos_i(7666) := b"1111111111111111_1111111111111111_1100000000011001_0010011001000000"; -- -0.24961625039577484
	pesos_i(7667) := b"0000000000000000_0000000000000000_0011011010110001_0011010000000000"; -- 0.21364140510559082
	pesos_i(7668) := b"1111111111111111_1111111111111111_1100010000111010_1010110100000000"; -- -0.23347967863082886
	pesos_i(7669) := b"0000000000000000_0000000000000000_0001011110001111_0111000110100000"; -- 0.0920325294137001
	pesos_i(7670) := b"1111111111111111_1111111111111111_0110100100101011_0101010000000000"; -- -0.5891826152801514
	pesos_i(7671) := b"0000000000000000_0000000000000000_0101100010000101_1100111110000000"; -- 0.3457917869091034
	pesos_i(7672) := b"1111111111111111_1111111111111111_0011111110010110_1000001100000000"; -- -0.7516096234321594
	pesos_i(7673) := b"0000000000000000_0000000000000000_0011011010100001_0011110011000000"; -- 0.2133977860212326
	pesos_i(7674) := b"1111111111111111_1111111111111111_1010100110000100_1100000000000000"; -- -0.3378181457519531
	pesos_i(7675) := b"0000000000000000_0000000000000000_0110001110100000_0001101100000000"; -- 0.38916176557540894
	pesos_i(7676) := b"1111111111111111_1111111111111111_1101000000001100_1010011011000000"; -- -0.1873069554567337
	pesos_i(7677) := b"1111111111111111_1111111111111111_1101010011010000_0100010110000000"; -- -0.1686970293521881
	pesos_i(7678) := b"0000000000000000_0000000000000000_0101100010010111_1111000100000000"; -- 0.34606844186782837
	pesos_i(7679) := b"0000000000000000_0000000000000000_0010100110001000_1011101001000000"; -- 0.16224254667758942
	pesos_i(7680) := b"1111111111111111_1111111111111111_1110011101110011_1101110110100000"; -- -0.09588827937841415
	pesos_i(7681) := b"0000000000000000_0000000000000000_1110101010011101_0100111100000000"; -- 0.9164628386497498
	pesos_i(7682) := b"0000000000000000_0000000000000000_0001000010001101_0110110101000000"; -- 0.06465800106525421
	pesos_i(7683) := b"0000000000000000_0000000000000000_0111101001011100_0010110110000000"; -- 0.4779690206050873
	pesos_i(7684) := b"1111111111111111_1111111111111111_1101011001100010_1010000111000000"; -- -0.16255749762058258
	pesos_i(7685) := b"0000000000000000_0000000000000000_0011111101111101_0000001011000000"; -- 0.24800126254558563
	pesos_i(7686) := b"0000000000000000_0000000000000000_0000010110001011_0011000111110000"; -- 0.02165519818663597
	pesos_i(7687) := b"1111111111111111_1111111111111111_1111000111101010_0100110110010000"; -- -0.05501857027411461
	pesos_i(7688) := b"0000000000000000_0000000000000000_0001001011101101_0100000000000000"; -- 0.07393264770507812
	pesos_i(7689) := b"0000000000000000_0000000000000000_0011101011011111_1001001110000000"; -- 0.22997400164604187
	pesos_i(7690) := b"0000000000000000_0000000000000000_1001010100100111_0001010000000000"; -- 0.582627534866333
	pesos_i(7691) := b"0000000000000000_0000000000000000_0100110110001111_0010100110000000"; -- 0.3029657304286957
	pesos_i(7692) := b"1111111111111111_1111111111111111_1110111100000010_1000111100000000"; -- -0.06636720895767212
	pesos_i(7693) := b"1111111111111111_1111111111111111_0010101111011110_1001100100000000"; -- -0.8286346793174744
	pesos_i(7694) := b"1111111111111111_1111111111111111_0000010101011101_1111001100000000"; -- -0.9790351986885071
	pesos_i(7695) := b"0000000000000000_0000000000000000_0001101011111111_0111110011100000"; -- 0.10546093434095383
	pesos_i(7696) := b"0000000000000000_0000000000000000_0001101101010001_1011100100100000"; -- 0.10671574622392654
	pesos_i(7697) := b"1111111111111111_1111111111111111_1110101000011110_0110010110000000"; -- -0.0854736864566803
	pesos_i(7698) := b"0000000000000000_0000000000000000_0001110010010001_0010001010100000"; -- 0.11158958822488785
	pesos_i(7699) := b"1111111111111111_1111111111111111_1001111011000101_1100101010000000"; -- -0.3797944486141205
	pesos_i(7700) := b"0000000000000000_0000000000000000_0001010001110111_0101100111100000"; -- 0.07994615286588669
	pesos_i(7701) := b"1111111111111111_1111111111111111_1100100001010001_1000110111000000"; -- -0.2175055891275406
	pesos_i(7702) := b"0000000000000000_0000000000000000_0110001100010111_0111001110000000"; -- 0.38707658648490906
	pesos_i(7703) := b"1111111111111111_1111111111111111_1110110010000011_1011010100100000"; -- -0.07611530274152756
	pesos_i(7704) := b"1111111111111111_1111111111111111_1111110101100000_0011011011100100"; -- -0.010250634513795376
	pesos_i(7705) := b"0000000000000000_0000000000000000_0101101100101101_0101110110000000"; -- 0.356160968542099
	pesos_i(7706) := b"1111111111111111_1111111111111111_1101111010010001_1000010101000000"; -- -0.13059203326702118
	pesos_i(7707) := b"1111111111111111_1111111111111111_1101010100011110_0010011010000000"; -- -0.16750869154930115
	pesos_i(7708) := b"0000000000000000_0000000000000000_0000000011011011_1100100111111101"; -- 0.003353714244440198
	pesos_i(7709) := b"1111111111111111_1111111111111111_1111110110100010_0111100100011100"; -- -0.009239607490599155
	pesos_i(7710) := b"0000000000000000_0000000000000000_1010011101010000_0110110100000000"; -- 0.6535709500312805
	pesos_i(7711) := b"0000000000000000_0000000000000000_0100011001101110_1101110100000000"; -- 0.27512913942337036
	pesos_i(7712) := b"1111111111111111_1111111111111111_1000000111001011_0111011110000000"; -- -0.49298909306526184
	pesos_i(7713) := b"1111111111111111_1111111111111111_1001000100010110_0001001000000000"; -- -0.43325698375701904
	pesos_i(7714) := b"0000000000000000_0000000000000000_0000010011100010_1000000010010000"; -- 0.019081149250268936
	pesos_i(7715) := b"0000000000000000_0000000000000000_0101010111000000_0000011100000000"; -- 0.3349613547325134
	pesos_i(7716) := b"1111111111111111_1111111111111111_1011000100011011_0111001110000000"; -- -0.30817487835884094
	pesos_i(7717) := b"0000000000000000_0000000000000000_0001010101011100_1110101111000000"; -- 0.0834491103887558
	pesos_i(7718) := b"1111111111111111_1111111111111111_1111010010001100_0010100111000000"; -- -0.04473628103733063
	pesos_i(7719) := b"0000000000000000_0000000000000000_1000000010001000_0001110000000000"; -- 0.5020768642425537
	pesos_i(7720) := b"0000000000000000_0000000000000000_0010000100110011_0111000101000000"; -- 0.1296911984682083
	pesos_i(7721) := b"1111111111111111_1111111111111111_1100101000111011_1010011110000000"; -- -0.21002724766731262
	pesos_i(7722) := b"1111111111111111_1111111111111111_1010000011110011_0110010010000000"; -- -0.3712861239910126
	pesos_i(7723) := b"0000000000000000_0000000000000000_0001011010101110_0101010101100000"; -- 0.0885976180434227
	pesos_i(7724) := b"0000000000000000_0000000000000000_0001111000110111_0010100001000000"; -- 0.11802913248538971
	pesos_i(7725) := b"0000000000000000_0000000000000000_0000110111010010_1011000100010000"; -- 0.05399614945054054
	pesos_i(7726) := b"0000000000000000_0000000000000000_0010010110010000_0111110101000000"; -- 0.14673598110675812
	pesos_i(7727) := b"0000000000000000_0000000000000000_1001111000010010_1011011100000000"; -- 0.6174730658531189
	pesos_i(7728) := b"1111111111111111_1111111111111111_1111111000010101_0011101011011110"; -- -0.007488556671887636
	pesos_i(7729) := b"1111111111111111_1111111111111111_0111101001000011_0110101000000000"; -- -0.5224088430404663
	pesos_i(7730) := b"0000000000000000_0000000000000000_0001000000111001_0001101110000000"; -- 0.06337139010429382
	pesos_i(7731) := b"0000000000000000_0000000000000000_0110000100110000_0001001010000000"; -- 0.37963977456092834
	pesos_i(7732) := b"0000000000000000_0000000000000000_1000100101011001_1001000100000000"; -- 0.5365229249000549
	pesos_i(7733) := b"1111111111111111_1111111111111111_1110110111111101_0011101001000000"; -- -0.07035480439662933
	pesos_i(7734) := b"0000000000000000_0000000000000000_0000100001010100_1110110100110000"; -- 0.03254587575793266
	pesos_i(7735) := b"0000000000000000_0000000000000000_1011000010101010_0000100000000000"; -- 0.6900944709777832
	pesos_i(7736) := b"0000000000000000_0000000000000000_0100011100010010_1010111000000000"; -- 0.2776287794113159
	pesos_i(7737) := b"0000000000000000_0000000000000000_1000011111000100_0101011000000000"; -- 0.5303395986557007
	pesos_i(7738) := b"0000000000000000_0000000000000000_0100101110001101_0010101110000000"; -- 0.29512283205986023
	pesos_i(7739) := b"0000000000000000_0000000000000000_0100101010101000_1111111110000000"; -- 0.2916412055492401
	pesos_i(7740) := b"0000000000000000_0000000000000000_0001011101111101_0011010011100000"; -- 0.091754250228405
	pesos_i(7741) := b"1111111111111111_1111111111111111_1000110000010100_1001100100000000"; -- -0.45281070470809937
	pesos_i(7742) := b"0000000000000000_0000000000000000_0111101110011100_1111000010000000"; -- 0.4828634560108185
	pesos_i(7743) := b"1111111111111111_1111111111111111_0011001100010011_1111101100000000"; -- -0.8004763722419739
	pesos_i(7744) := b"0000000000000000_0000000000000000_0000010100001000_0110101100001000"; -- 0.019659699872136116
	pesos_i(7745) := b"1111111111111111_1111111111111111_1101011000111011_0001110001000000"; -- -0.1631605476140976
	pesos_i(7746) := b"0000000000000000_0000000000000000_0011001100011110_0011000011000000"; -- 0.1996794193983078
	pesos_i(7747) := b"0000000000000000_0000000000000000_0010100001010110_1001001011000000"; -- 0.1575710028409958
	pesos_i(7748) := b"0000000000000000_0000000000000000_0001100110010001_0110001110000000"; -- 0.09987470507621765
	pesos_i(7749) := b"1111111111111111_1111111111111111_1100100111010101_1001001000000000"; -- -0.2115849256515503
	pesos_i(7750) := b"0000000000000000_0000000000000000_0011100010011110_0101000011000000"; -- 0.2211657017469406
	pesos_i(7751) := b"1111111111111111_1111111111111111_1101001110110101_1100111010000000"; -- -0.17300710082054138
	pesos_i(7752) := b"1111111111111111_1111111111111111_1000001101111011_0111100110000000"; -- -0.4863971769809723
	pesos_i(7753) := b"0000000000000000_0000000000000000_1010010011111001_0000001000000000"; -- 0.644424557685852
	pesos_i(7754) := b"1111111111111111_1111111111111111_1110111100100101_1101101011000000"; -- -0.06582863628864288
	pesos_i(7755) := b"1111111111111111_1111111111111111_1000011100100001_0000110000000000"; -- -0.4721519947052002
	pesos_i(7756) := b"0000000000000000_0000000000000000_0001001101110011_1001001111100000"; -- 0.07598232477903366
	pesos_i(7757) := b"0000000000000000_0000000000000000_0011101011011001_1001111101000000"; -- 0.22988314926624298
	pesos_i(7758) := b"1111111111111111_1111111111111111_1000101001110111_0111111000000000"; -- -0.4591141939163208
	pesos_i(7759) := b"1111111111111111_1111111111111111_1100101110111001_1101111010000000"; -- -0.20419511198997498
	pesos_i(7760) := b"1111111111111111_1111111111111111_1111000111001101_0011110001000000"; -- -0.05546210706233978
	pesos_i(7761) := b"0000000000000000_0000000000000000_0100011100001000_0001011000000000"; -- 0.27746713161468506
	pesos_i(7762) := b"1111111111111111_1111111111111111_0110110101110110_0010101100000000"; -- -0.5724156498908997
	pesos_i(7763) := b"1111111111111111_1111111111111111_0101111110000001_1111110100000000"; -- -0.6269227862358093
	pesos_i(7764) := b"0000000000000000_0000000000000000_0101111010101011_1111101100000000"; -- 0.3698117136955261
	pesos_i(7765) := b"0000000000000000_0000000000000000_1010100011111000_0100111000000000"; -- 0.6600388288497925
	pesos_i(7766) := b"1111111111111111_1111111111111111_1101010000011001_0101100000000000"; -- -0.17148828506469727
	pesos_i(7767) := b"0000000000000000_0000000000000000_0010010000101010_1011101010000000"; -- 0.1412769854068756
	pesos_i(7768) := b"0000000000000000_0000000000000000_0110000000001100_0100111110000000"; -- 0.37518784403800964
	pesos_i(7769) := b"1111111111111111_1111111111111111_0110101110000010_0100100100000000"; -- -0.5800432562828064
	pesos_i(7770) := b"1111111111111111_1111111111111111_1000111011001100_1111101010000000"; -- -0.44218477606773376
	pesos_i(7771) := b"0000000000000000_0000000000000000_0010100111101110_0011000011000000"; -- 0.1637907475233078
	pesos_i(7772) := b"0000000000000000_0000000000000000_0010101000111100_0010100001000000"; -- 0.1649804264307022
	pesos_i(7773) := b"0000000000000000_0000000000000000_0101111001001111_1011011010000000"; -- 0.368403822183609
	pesos_i(7774) := b"0000000000000000_0000000000000000_0010110110011000_1111010010000000"; -- 0.17811515927314758
	pesos_i(7775) := b"1111111111111111_1111111111111111_1010101111010111_0011010000000000"; -- -0.3287475109100342
	pesos_i(7776) := b"0000000000000000_0000000000000000_0110100001001111_0011000110000000"; -- 0.4074583947658539
	pesos_i(7777) := b"0000000000000000_0000000000000000_0000101010011100_0001011001000000"; -- 0.04144419729709625
	pesos_i(7778) := b"0000000000000000_0000000000000000_0101110000010000_1111110100000000"; -- 0.3596342206001282
	pesos_i(7779) := b"0000000000000000_0000000000000000_0001000000001111_1000111011000000"; -- 0.06273739039897919
	pesos_i(7780) := b"0000000000000000_0000000000000000_0001100000101011_1100100010100000"; -- 0.09441808611154556
	pesos_i(7781) := b"1111111111111111_1111111111111111_1000111100100011_0000010000000000"; -- -0.4408719539642334
	pesos_i(7782) := b"1111111111111111_1111111111111111_1101101000100010_1110110101000000"; -- -0.14790455996990204
	pesos_i(7783) := b"1111111111111111_1111111111111111_1000110101000111_1011011000000000"; -- -0.4481245279312134
	pesos_i(7784) := b"0000000000000000_0000000000000000_0000100011101100_1110101111000000"; -- 0.0348651260137558
	pesos_i(7785) := b"1111111111111111_1111111111111111_1111101110000011_0100010101011000"; -- -0.017528215423226357
	pesos_i(7786) := b"0000000000000000_0000000000000000_1001011000010100_0101011100000000"; -- 0.5862478613853455
	pesos_i(7787) := b"1111111111111111_1111111111111111_1000100111011010_0011101000000000"; -- -0.461513876914978
	pesos_i(7788) := b"1111111111111111_1111111111111111_1101011110111110_0111011000000000"; -- -0.1572500467300415
	pesos_i(7789) := b"0000000000000000_0000000000000000_0010010111010001_0100111011000000"; -- 0.14772503077983856
	pesos_i(7790) := b"1111111111111111_1111111111111111_1100011100011100_1000000101000000"; -- -0.22222130000591278
	pesos_i(7791) := b"0000000000000000_0000000000000000_0010001110001010_0011011101000000"; -- 0.13882775604724884
	pesos_i(7792) := b"1111111111111111_1111111111111111_1001011111111110_0101011100000000"; -- -0.40627533197402954
	pesos_i(7793) := b"0000000000000000_0000000000000000_0010011011100101_1000011001000000"; -- 0.1519397646188736
	pesos_i(7794) := b"1111111111111111_1111111111111111_1010010000101101_0101010100000000"; -- -0.3586832880973816
	pesos_i(7795) := b"0000000000000000_0000000000000000_0000111010001100_1011011101000000"; -- 0.05683465301990509
	pesos_i(7796) := b"0000000000000000_0000000000000000_0011110010111100_1111100011000000"; -- 0.23725847899913788
	pesos_i(7797) := b"0000000000000000_0000000000000000_0001100001100110_1011001101000000"; -- 0.09531708061695099
	pesos_i(7798) := b"1111111111111111_1111111111111111_0111110011100011_0110011000000000"; -- -0.5121551752090454
	pesos_i(7799) := b"1111111111111111_1111111111111111_1110110101001000_1000110001000000"; -- -0.07311175763607025
	pesos_i(7800) := b"1111111111111111_1111111111111111_0111000001011110_1110011100000000"; -- -0.5610519051551819
	pesos_i(7801) := b"0000000000000000_0000000000000000_0001000100001011_0010110101000000"; -- 0.06657679378986359
	pesos_i(7802) := b"1111111111111111_1111111111111111_1011100110000101_0111001110000000"; -- -0.27530744671821594
	pesos_i(7803) := b"0000000000000000_0000000000000000_0101000010011100_0010110010000000"; -- 0.3148830235004425
	pesos_i(7804) := b"1111111111111111_1111111111111111_1011111010101001_1001111110000000"; -- -0.2552242577075958
	pesos_i(7805) := b"1111111111111111_1111111111111111_1000010111010101_1100101100000000"; -- -0.4772065281867981
	pesos_i(7806) := b"1111111111111111_1111111111111111_1111111111111110_0111111101110110"; -- -2.2920314222574234e-05
	pesos_i(7807) := b"1111111111111111_1111111111111111_1111100011111010_1101010000001000"; -- -0.027422664687037468
	pesos_i(7808) := b"1111111111111111_1111111111111111_0101110110010000_0101010000000000"; -- -0.6345164775848389
	pesos_i(7809) := b"0000000000000000_0000000000000000_0110010011110111_1111101010000000"; -- 0.39440885186195374
	pesos_i(7810) := b"0000000000000000_0000000000000000_0010110101000111_1010111110000000"; -- 0.17687508463859558
	pesos_i(7811) := b"0000000000000000_0000000000000000_0011010010011010_1111100001000000"; -- 0.2054896503686905
	pesos_i(7812) := b"1111111111111111_1111111111111111_1101101101000011_0101110110000000"; -- -0.143503338098526
	pesos_i(7813) := b"0000000000000000_0000000000000000_0010100010010010_1111001100000000"; -- 0.15849226713180542
	pesos_i(7814) := b"1111111111111111_1111111111111111_1101110000010110_0101101101000000"; -- -0.14028386771678925
	pesos_i(7815) := b"0000000000000000_0000000000000000_0000111101111100_1100111010010000"; -- 0.06049815192818642
	pesos_i(7816) := b"0000000000000000_0000000000000000_0000000000000111_1110011110101110"; -- 0.00012062069436069578
	pesos_i(7817) := b"1111111111111111_1111111111111111_1110100001110001_1100001011000000"; -- -0.09201414883136749
	pesos_i(7818) := b"0000000000000000_0000000000000000_0010010110111001_0110000000000000"; -- 0.14735984802246094
	pesos_i(7819) := b"0000000000000000_0000000000000000_0000100010111110_1100000010100000"; -- 0.03416065126657486
	pesos_i(7820) := b"1111111111111111_1111111111111111_1111011101010000_1111001000000000"; -- -0.033921122550964355
	pesos_i(7821) := b"1111111111111111_1111111111111111_1000000010010001_1110011110000000"; -- -0.497773677110672
	pesos_i(7822) := b"1111111111111111_1111111111111111_0011111111001110_0110111000000000"; -- -0.7507563829421997
	pesos_i(7823) := b"1111111111111111_1111111111111111_1111101001000001_1110100100001000"; -- -0.022431788966059685
	pesos_i(7824) := b"0000000000000000_0000000000000000_0101001000110000_1000110110000000"; -- 0.3210533559322357
	pesos_i(7825) := b"1111111111111111_1111111111111111_1001101001111110_0111100000000000"; -- -0.39650774002075195
	pesos_i(7826) := b"0000000000000000_0000000000000000_0000101000110101_0011100101000000"; -- 0.03987462818622589
	pesos_i(7827) := b"1111111111111111_1111111111111111_0111100001100110_1010010100000000"; -- -0.5296837687492371
	pesos_i(7828) := b"1111111111111111_1111111111111111_1111011101110111_0001100101010000"; -- -0.03333894535899162
	pesos_i(7829) := b"0000000000000000_0000000000000000_0000110111111001_0000111000100000"; -- 0.05458153039216995
	pesos_i(7830) := b"0000000000000000_0000000000000000_0001101110100110_0101010010100000"; -- 0.10800675302743912
	pesos_i(7831) := b"0000000000000000_0000000000000000_0010011000101100_1100010100000000"; -- 0.14912062883377075
	pesos_i(7832) := b"0000000000000000_0000000000000000_0010001000101011_0101010011000000"; -- 0.13347367942333221
	pesos_i(7833) := b"0000000000000000_0000000000000000_0100110011111110_1000111010000000"; -- 0.3007592260837555
	pesos_i(7834) := b"1111111111111111_1111111111111111_1100101101111111_1000010110000000"; -- -0.20508542656898499
	pesos_i(7835) := b"1111111111111111_1111111111111111_0101100100011011_0011101000000000"; -- -0.6519283056259155
	pesos_i(7836) := b"0000000000000000_0000000000000000_0000101001111010_1101000100010000"; -- 0.040936533361673355
	pesos_i(7837) := b"0000000000000000_0000000000000000_0000100101001100_0100010110110000"; -- 0.036320071667432785
	pesos_i(7838) := b"0000000000000000_0000000000000000_0001110101011100_0010111110100000"; -- 0.11468789726495743
	pesos_i(7839) := b"0000000000000000_0000000000000000_0001101100011100_0111011011100000"; -- 0.10590308159589767
	pesos_i(7840) := b"1111111111111111_1111111111111111_0111110100001011_0011101100000000"; -- -0.5115473866462708
	pesos_i(7841) := b"0000000000000000_0000000000000000_0000001011101100_0100101110111100"; -- 0.011418088339269161
	pesos_i(7842) := b"1111111111111111_1111111111111111_1011101001011100_0111010010000000"; -- -0.27202674746513367
	pesos_i(7843) := b"0000000000000000_0000000000000000_0001110111000100_1011101101000000"; -- 0.11628313362598419
	pesos_i(7844) := b"1111111111111111_1111111111111111_1011100111101001_1010001010000000"; -- -0.2737787663936615
	pesos_i(7845) := b"1111111111111111_1111111111111111_1100111110100100_1010000111000000"; -- -0.18889416754245758
	pesos_i(7846) := b"1111111111111111_1111111111111111_1001101101011111_1010100100000000"; -- -0.39307159185409546
	pesos_i(7847) := b"0000000000000000_0000000000000000_0011100001101101_1000111100000000"; -- 0.22042173147201538
	pesos_i(7848) := b"1111111111111111_1111111111111111_1110001111101101_1001100111000000"; -- -0.10965575277805328
	pesos_i(7849) := b"0000000000000000_0000000000000000_0001001000000101_1010111101000000"; -- 0.07039923965930939
	pesos_i(7850) := b"1111111111111111_1111111111111111_0110111111111011_1000001100000000"; -- -0.5625684857368469
	pesos_i(7851) := b"0000000000000000_0000000000000000_0010011011001001_1011011000000000"; -- 0.15151536464691162
	pesos_i(7852) := b"0000000000000000_0000000000000000_0011000010001100_0000011111000000"; -- 0.189636692404747
	pesos_i(7853) := b"1111111111111111_1111111111111111_1111000000111111_1011011001010000"; -- -0.06152782961726189
	pesos_i(7854) := b"0000000000000000_0000000000000000_1000001101100111_1110011000000000"; -- 0.5133041143417358
	pesos_i(7855) := b"0000000000000000_0000000000000000_0110000110010101_0010011010000000"; -- 0.38118210434913635
	pesos_i(7856) := b"1111111111111111_1111111111111111_1100110010001000_1100111011000000"; -- -0.2010374814271927
	pesos_i(7857) := b"1111111111111111_1111111111111111_1000111011101011_1010011000000000"; -- -0.4417167901992798
	pesos_i(7858) := b"1111111111111111_1111111111111111_1101101010010000_0110010111000000"; -- -0.1462341696023941
	pesos_i(7859) := b"0000000000000000_0000000000000000_0101001100110001_0110001110000000"; -- 0.32497236132621765
	pesos_i(7860) := b"0000000000000000_0000000000000000_0101011101000010_1011110010000000"; -- 0.34086206555366516
	pesos_i(7861) := b"1111111111111111_1111111111111111_1110010010110110_1101011110100000"; -- -0.1065850481390953
	pesos_i(7862) := b"1111111111111111_1111111111111111_1101000111001111_1100011100000000"; -- -0.1804233193397522
	pesos_i(7863) := b"0000000000000000_0000000000000000_1000010111110010_0110000100000000"; -- 0.5232296586036682
	pesos_i(7864) := b"0000000000000000_0000000000000000_0001010110011010_0100011100000000"; -- 0.08438533544540405
	pesos_i(7865) := b"0000000000000000_0000000000000000_0011001100011010_0011111110000000"; -- 0.19961926341056824
	pesos_i(7866) := b"0000000000000000_0000000000000000_0001011101001000_0010011110100000"; -- 0.09094474464654922
	pesos_i(7867) := b"1111111111111111_1111111111111111_1010111011010011_0100001100000000"; -- -0.31708890199661255
	pesos_i(7868) := b"1111111111111111_1111111111111111_1111110000010100_0110001101101000"; -- -0.015313899144530296
	pesos_i(7869) := b"0000000000000000_0000000000000000_0001100010111001_0101100010100000"; -- 0.09657815843820572
	pesos_i(7870) := b"1111111111111111_1111111111111111_1110101001000100_0111111100000000"; -- -0.08489233255386353
	pesos_i(7871) := b"1111111111111111_1111111111111111_0011010011000010_0011001100000000"; -- -0.7939117550849915
	pesos_i(7872) := b"1111111111111111_1111111111111111_1111011001111000_1100011100100000"; -- -0.0372195765376091
	pesos_i(7873) := b"1111111111111111_1111111111111111_1101100000000001_0001011110000000"; -- -0.15623334050178528
	pesos_i(7874) := b"0000000000000000_0000000000000000_0000101111000001_0100100101110000"; -- 0.04591807350516319
	pesos_i(7875) := b"0000000000000000_0000000000000000_0010000110100101_1001011111000000"; -- 0.13143299520015717
	pesos_i(7876) := b"0000000000000000_0000000000000000_0011101110100000_0000101110000000"; -- 0.23291084170341492
	pesos_i(7877) := b"1111111111111111_1111111111111111_1010001100100100_1001101000000000"; -- -0.3627227544784546
	pesos_i(7878) := b"1111111111111111_1111111111111111_1101000110101001_1101100010000000"; -- -0.18100211024284363
	pesos_i(7879) := b"0000000000000000_0000000000000000_0011000010000000_0101101000000000"; -- 0.18945848941802979
	pesos_i(7880) := b"1111111111111111_1111111111111111_1010100000110011_1100001110000000"; -- -0.3429601490497589
	pesos_i(7881) := b"0000000000000000_0000000000000000_1000000000001000_1101101100000000"; -- 0.5001351237297058
	pesos_i(7882) := b"0000000000000000_0000000000000000_0000101010001110_1000011100010000"; -- 0.041237298399209976
	pesos_i(7883) := b"1111111111111111_1111111111111111_0111001010011100_1011001100000000"; -- -0.5522964596748352
	pesos_i(7884) := b"1111111111111111_1111111111111111_1110000010111011_0001000110100000"; -- -0.12214555591344833
	pesos_i(7885) := b"0000000000000000_0000000000000000_0101100110111111_0100011100000000"; -- 0.35057491064071655
	pesos_i(7886) := b"1111111111111111_1111111111111111_1001000001111000_0110110100000000"; -- -0.4356624484062195
	pesos_i(7887) := b"1111111111111111_1111111111111111_1001011100110101_1101111010000000"; -- -0.409334272146225
	pesos_i(7888) := b"0000000000000000_0000000000000000_0010110010011000_0011100101000000"; -- 0.1741977483034134
	pesos_i(7889) := b"0000000000000000_0000000000000000_0010110010110010_1000110101000000"; -- 0.17459948360919952
	pesos_i(7890) := b"1111111111111111_1111111111111111_0110110100010001_0011000000000000"; -- -0.5739564895629883
	pesos_i(7891) := b"1111111111111111_1111111111111111_1100110000011101_1111010101000000"; -- -0.20266787707805634
	pesos_i(7892) := b"0000000000000000_0000000000000000_0010100000000101_1111001101000000"; -- 0.1563407927751541
	pesos_i(7893) := b"0000000000000000_0000000000000000_0100111101111100_1111000010000000"; -- 0.3105001747608185
	pesos_i(7894) := b"0000000000000000_0000000000000000_0001001111000001_0100101011000000"; -- 0.07716815173625946
	pesos_i(7895) := b"0000000000000000_0000000000000000_0000010101101110_1110101101110000"; -- 0.021223749965429306
	pesos_i(7896) := b"0000000000000000_0000000000000000_0011000010101011_1000000101000000"; -- 0.19011695683002472
	pesos_i(7897) := b"1111111111111111_1111111111111111_0111100010011001_0110101000000000"; -- -0.5289090871810913
	pesos_i(7898) := b"0000000000000000_0000000000000000_0000110110101010_1010010010010000"; -- 0.05338505282998085
	pesos_i(7899) := b"1111111111111111_1111111111111111_1101010000011000_1111101000000000"; -- -0.17149388790130615
	pesos_i(7900) := b"1111111111111111_1111111111111111_1001000011100011_0100101100000000"; -- -0.43403178453445435
	pesos_i(7901) := b"0000000000000000_0000000000000000_0110000100010011_1001111000000000"; -- 0.379205584526062
	pesos_i(7902) := b"0000000000000000_0000000000000000_0011011101001010_0101100010000000"; -- 0.21597817540168762
	pesos_i(7903) := b"0000000000000000_0000000000000000_0001000110111110_1100010101100000"; -- 0.06931718438863754
	pesos_i(7904) := b"0000000000000000_0000000000000000_0100010000000001_1101101100000000"; -- 0.2656533122062683
	pesos_i(7905) := b"1111111111111111_1111111111111111_1111110001010011_1101111111000000"; -- -0.014345183968544006
	pesos_i(7906) := b"0000000000000000_0000000000000000_0110101010101110_0001001110000000"; -- 0.4167186915874481
	pesos_i(7907) := b"1111111111111111_1111111111111111_1101111101100111_1110111111000000"; -- -0.1273203045129776
	pesos_i(7908) := b"0000000000000000_0000000000000000_0000010011110110_0010101000000000"; -- 0.019381165504455566
	pesos_i(7909) := b"1111111111111111_1111111111111111_1111010000001011_1111011110010000"; -- -0.04669239744544029
	pesos_i(7910) := b"1111111111111111_1111111111111111_1011000100001101_1001101010000000"; -- -0.3083861768245697
	pesos_i(7911) := b"1111111111111111_1111111111111111_0110000111100100_1110000100000000"; -- -0.6176013350486755
	pesos_i(7912) := b"0000000000000000_0000000000000000_0100011101001001_0001011010000000"; -- 0.27845898270606995
	pesos_i(7913) := b"0000000000000000_0000000000000000_0000001101111010_1010110110001000"; -- 0.01359066553413868
	pesos_i(7914) := b"0000000000000000_0000000000000000_0011100011111011_1010010010000000"; -- 0.22258976101875305
	pesos_i(7915) := b"1111111111111111_1111111111111111_1011101111001100_1000111010000000"; -- -0.2664099633693695
	pesos_i(7916) := b"1111111111111111_1111111111111111_1110111100010001_1110111101000000"; -- -0.06613259017467499
	pesos_i(7917) := b"0000000000000000_0000000000000000_0110010011100100_0011101100000000"; -- 0.39410752058029175
	pesos_i(7918) := b"1111111111111111_1111111111111111_0100001111110111_1101110000000000"; -- -0.7344992160797119
	pesos_i(7919) := b"0000000000000000_0000000000000000_0001000101110100_0010010101000000"; -- 0.06817848980426788
	pesos_i(7920) := b"1111111111111111_1111111111111111_1100110100010101_1011001011000000"; -- -0.1988876610994339
	pesos_i(7921) := b"0000000000000000_0000000000000000_0001011001011110_0010000000100000"; -- 0.08737374097108841
	pesos_i(7922) := b"1111111111111111_1111111111111111_0111000000001010_0111011000000000"; -- -0.5623403787612915
	pesos_i(7923) := b"0000000000000000_0000000000000000_0011011101101000_1011110110000000"; -- 0.21644195914268494
	pesos_i(7924) := b"0000000000000000_0000000000000000_0000101000010001_1001001111100000"; -- 0.03933071345090866
	pesos_i(7925) := b"0000000000000000_0000000000000000_0010010000011100_1101010111000000"; -- 0.14106498658657074
	pesos_i(7926) := b"0000000000000000_0000000000000000_0000000100100000_0000011101101010"; -- 0.004394973162561655
	pesos_i(7927) := b"0000000000000000_0000000000000000_0000000111001111_0000001001001000"; -- 0.007064955309033394
	pesos_i(7928) := b"1111111111111111_1111111111111111_1011000110010100_1101111110000000"; -- -0.3063221275806427
	pesos_i(7929) := b"1111111111111111_1111111111111111_1101101111111001_0000000101000000"; -- -0.14073173701763153
	pesos_i(7930) := b"1111111111111111_1111111111111111_1100011001000111_1110101000000000"; -- -0.22546517848968506
	pesos_i(7931) := b"0000000000000000_0000000000000000_0011000110110001_0111111111000000"; -- 0.19411467015743256
	pesos_i(7932) := b"1111111111111111_1111111111111111_1101011011110110_0010010100000000"; -- -0.1603066325187683
	pesos_i(7933) := b"0000000000000000_0000000000000000_0001001110010100_0011010110000000"; -- 0.07648023962974548
	pesos_i(7934) := b"0000000000000000_0000000000000000_0000001000001011_1101001100111000"; -- 0.007992936298251152
	pesos_i(7935) := b"0000000000000000_0000000000000000_0101101010011010_0011011010000000"; -- 0.35391560196876526
	pesos_i(7936) := b"1111111111111111_1111111111111111_1010000101100100_0001001000000000"; -- -0.36956679821014404
	pesos_i(7937) := b"0000000000000000_0000000000000000_0010011011000000_0110101001000000"; -- 0.15137352049350739
	pesos_i(7938) := b"1111111111111111_1111111111111111_1100101011010000_0010000110000000"; -- -0.20776167511940002
	pesos_i(7939) := b"0000000000000000_0000000000000000_0001001000001010_1011011100000000"; -- 0.0704759955406189
	pesos_i(7940) := b"1111111111111111_1111111111111111_1110101110011011_1110011110000000"; -- -0.079652339220047
	pesos_i(7941) := b"1111111111111111_1111111111111111_1100101001001001_1011101110000000"; -- -0.20981243252754211
	pesos_i(7942) := b"1111111111111111_1111111111111111_1111100101110110_0011010101011000"; -- -0.025540033355355263
	pesos_i(7943) := b"1111111111111111_1111111111111111_1111111001110100_1110011110101010"; -- -0.006028672214597464
	pesos_i(7944) := b"1111111111111111_1111111111111111_1110010101111000_0001010111100000"; -- -0.10363639146089554
	pesos_i(7945) := b"0000000000000000_0000000000000000_0011001010101011_0011111111000000"; -- 0.19792555272579193
	pesos_i(7946) := b"1111111111111111_1111111111111111_1101010010110000_0000100000000000"; -- -0.1691889762878418
	pesos_i(7947) := b"1111111111111111_1111111111111111_1101001001001110_0000010110000000"; -- -0.17849698662757874
	pesos_i(7948) := b"1111111111111111_1111111111111111_1111110110101100_1001000011011100"; -- -0.00908560398966074
	pesos_i(7949) := b"1111111111111111_1111111111111111_1100000011101011_1111111101000000"; -- -0.24639897048473358
	pesos_i(7950) := b"1111111111111111_1111111111111111_1101110110001100_0010100110000000"; -- -0.13458004593849182
	pesos_i(7951) := b"1111111111111111_1111111111111111_1110000011100000_1010101010100000"; -- -0.1215718612074852
	pesos_i(7952) := b"0000000000000000_0000000000000000_0010110100000011_0101000000000000"; -- 0.17583179473876953
	pesos_i(7953) := b"0000000000000000_0000000000000000_0001000001100000_0000100010100000"; -- 0.06396535784006119
	pesos_i(7954) := b"1111111111111111_1111111111111111_1111111111110010_0000100011010100"; -- -0.0002130968205165118
	pesos_i(7955) := b"1111111111111111_1111111111111111_1110110101011010_1001011110100000"; -- -0.07283642143011093
	pesos_i(7956) := b"0000000000000000_0000000000000000_0001001111100111_0001011111100000"; -- 0.07774495333433151
	pesos_i(7957) := b"0000000000000000_0000000000000000_0000010010110010_0001101100100000"; -- 0.018342681229114532
	pesos_i(7958) := b"1111111111111111_1111111111111111_1111101100110100_1100111110001000"; -- -0.018725423142313957
	pesos_i(7959) := b"0000000000000000_0000000000000000_0000101111011100_1101011111010000"; -- 0.04633854702115059
	pesos_i(7960) := b"1111111111111111_1111111111111111_1111011101000001_1110001011110000"; -- -0.034150902181863785
	pesos_i(7961) := b"0000000000000000_0000000000000000_0001111011010110_1111011001000000"; -- 0.12046755850315094
	pesos_i(7962) := b"1111111111111111_1111111111111111_1110010101110100_1000001011100000"; -- -0.10369092971086502
	pesos_i(7963) := b"1111111111111111_1111111111111111_1001000111000011_1011110100000000"; -- -0.43060702085494995
	pesos_i(7964) := b"0000000000000000_0000000000000000_0011001011100010_1011100110000000"; -- 0.19877204298973083
	pesos_i(7965) := b"1111111111111111_1111111111111111_1110001010101001_0010010100100000"; -- -0.11460655182600021
	pesos_i(7966) := b"1111111111111111_1111111111111111_1110110000001011_1011010011000000"; -- -0.07794637978076935
	pesos_i(7967) := b"1111111111111111_1111111111111111_1111101110111111_1010110011111000"; -- -0.016606511548161507
	pesos_i(7968) := b"1111111111111111_1111111111111111_1110001110101001_1101110111000000"; -- -0.11068929731845856
	pesos_i(7969) := b"0000000000000000_0000000000000000_0000101100000101_0001001101100000"; -- 0.04304619878530502
	pesos_i(7970) := b"1111111111111111_1111111111111111_1101111001100111_0101011100000000"; -- -0.13123565912246704
	pesos_i(7971) := b"0000000000000000_0000000000000000_0000111010111100_1010010111000000"; -- 0.05756603181362152
	pesos_i(7972) := b"1111111111111111_1111111111111111_1101110101110001_0011101110000000"; -- -0.13499096035957336
	pesos_i(7973) := b"1111111111111111_1111111111111111_1110010110100110_1001101001100000"; -- -0.1029265895485878
	pesos_i(7974) := b"0000000000000000_0000000000000000_0000110000001011_1100101100110000"; -- 0.0470549575984478
	pesos_i(7975) := b"1111111111111111_1111111111111111_1111011100011100_1100111101000000"; -- -0.0347166508436203
	pesos_i(7976) := b"1111111111111111_1111111111111111_1111100011000111_0001010010000000"; -- -0.028212279081344604
	pesos_i(7977) := b"1111111111111111_1111111111111111_1110100010010011_0011100100100000"; -- -0.0915035530924797
	pesos_i(7978) := b"1111111111111111_1111111111111111_1001010111111010_1011110010000000"; -- -0.41414281725883484
	pesos_i(7979) := b"1111111111111111_1111111111111111_1100100110010000_1001010000000000"; -- -0.21263766288757324
	pesos_i(7980) := b"0000000000000000_0000000000000000_0011100100000111_1100011001000000"; -- 0.22277487814426422
	pesos_i(7981) := b"0000000000000000_0000000000000000_0000011110111000_1101111011000000"; -- 0.030164644122123718
	pesos_i(7982) := b"0000000000000000_0000000000000000_0010111011001101_0000010011000000"; -- 0.18281583487987518
	pesos_i(7983) := b"0000000000000000_0000000000000000_0000000000011000_0000011000010011"; -- 0.00036657298915088177
	pesos_i(7984) := b"1111111111111111_1111111111111111_1010111101100110_1110000000000000"; -- -0.3148365020751953
	pesos_i(7985) := b"1111111111111111_1111111111111111_1010010011100101_0101111110000000"; -- -0.35587504506111145
	pesos_i(7986) := b"1111111111111111_1111111111111111_1100110111101010_1110100000000000"; -- -0.1956343650817871
	pesos_i(7987) := b"0000000000000000_0000000000000000_0001101000100110_1111011000100000"; -- 0.10215700417757034
	pesos_i(7988) := b"0000000000000000_0000000000000000_0000110000100100_0000110011110000"; -- 0.04742508754134178
	pesos_i(7989) := b"1111111111111111_1111111111111111_1101011100111101_1010111010000000"; -- -0.1592150628566742
	pesos_i(7990) := b"1111111111111111_1111111111111111_1111001011100111_1000001101010000"; -- -0.05115489289164543
	pesos_i(7991) := b"0000000000000000_0000000000000000_0001101111101010_0000001000100000"; -- 0.10903943330049515
	pesos_i(7992) := b"0000000000000000_0000000000000000_0000110100010111_0100001001010000"; -- 0.05113615468144417
	pesos_i(7993) := b"0000000000000000_0000000000000000_0000101100011100_1101011110110000"; -- 0.04340885207056999
	pesos_i(7994) := b"1111111111111111_1111111111111111_1110101110100011_1100111011000000"; -- -0.07953174412250519
	pesos_i(7995) := b"1111111111111111_1111111111111111_1001011100101110_1110011110000000"; -- -0.4094405472278595
	pesos_i(7996) := b"1111111111111111_1111111111111111_1110101010101010_1111011100000000"; -- -0.08332878351211548
	pesos_i(7997) := b"0000000000000000_0000000000000000_0010110100100110_0111110101000000"; -- 0.17636854946613312
	pesos_i(7998) := b"1111111111111111_1111111111111111_1110010100110001_1011111111100000"; -- -0.10470963269472122
	pesos_i(7999) := b"1111111111111111_1111111111111111_1100011010000000_0100110000000000"; -- -0.22460484504699707
	pesos_i(8000) := b"0000000000000000_0000000000000000_0000000001100101_1000101110011000"; -- 0.0015494580147787929
	pesos_i(8001) := b"0000000000000000_0000000000000000_0000101110011110_1101110111010000"; -- 0.04539285972714424
	pesos_i(8002) := b"0000000000000000_0000000000000000_0000010001011100_0011100010011000"; -- 0.017032181844115257
	pesos_i(8003) := b"0000000000000000_0000000000000000_0010011110110000_1011101111000000"; -- 0.15504048764705658
	pesos_i(8004) := b"1111111111111111_1111111111111111_1110101010000011_0110110001000000"; -- -0.08393214643001556
	pesos_i(8005) := b"1111111111111111_1111111111111111_1110101011111011_1000110101000000"; -- -0.08209912478923798
	pesos_i(8006) := b"0000000000000000_0000000000000000_0000100010000100_0101111011000000"; -- 0.03326980769634247
	pesos_i(8007) := b"0000000000000000_0000000000000000_0001101010101110_0001100110100000"; -- 0.10421905666589737
	pesos_i(8008) := b"1111111111111111_1111111111111111_1100011100011001_0111100100000000"; -- -0.22226756811141968
	pesos_i(8009) := b"0000000000000000_0000000000000000_0100000010111010_0110110000000000"; -- 0.25284457206726074
	pesos_i(8010) := b"0000000000000000_0000000000000000_0001100100101001_0100001101100000"; -- 0.09828587621450424
	pesos_i(8011) := b"1111111111111111_1111111111111111_1110000010111110_0001100111000000"; -- -0.12209929525852203
	pesos_i(8012) := b"0000000000000000_0000000000000000_0000110010000000_1000111110100000"; -- 0.048836685717105865
	pesos_i(8013) := b"0000000000000000_0000000000000000_0000101011111000_1111111001110000"; -- 0.04286184534430504
	pesos_i(8014) := b"1111111111111111_1111111111111111_1010111000101111_0110111110000000"; -- -0.31958869099617004
	pesos_i(8015) := b"1111111111111111_1111111111111111_1111010111011100_1010110000110000"; -- -0.03960155323147774
	pesos_i(8016) := b"0000000000000000_0000000000000000_0000011000111111_1011111110111000"; -- 0.024410231038928032
	pesos_i(8017) := b"0000000000000000_0000000000000000_0011000110000010_0100000011000000"; -- 0.1933937519788742
	pesos_i(8018) := b"1111111111111111_1111111111111111_1111010100000011_1100010110110000"; -- -0.042911190539598465
	pesos_i(8019) := b"0000000000000000_0000000000000000_0000010000011101_1101101001000000"; -- 0.01608051359653473
	pesos_i(8020) := b"1111111111111111_1111111111111111_1111000010010011_1110111101000000"; -- -0.06024269759654999
	pesos_i(8021) := b"0000000000000000_0000000000000000_0000010010001000_1110100011001000"; -- 0.01771407015621662
	pesos_i(8022) := b"0000000000000000_0000000000000000_0001001000010110_0000010101000000"; -- 0.07064850628376007
	pesos_i(8023) := b"0000000000000000_0000000000000000_0011000000100111_0111110010000000"; -- 0.18810251355171204
	pesos_i(8024) := b"0000000000000000_0000000000000000_0000111010101000_0100011100100000"; -- 0.05725521594285965
	pesos_i(8025) := b"1111111111111111_1111111111111111_1100010111000111_1010100100000000"; -- -0.22742217779159546
	pesos_i(8026) := b"1111111111111111_1111111111111111_1110001010011101_0010110110000000"; -- -0.11478915810585022
	pesos_i(8027) := b"0000000000000000_0000000000000000_0000010111000110_1010000100110000"; -- 0.022562097758054733
	pesos_i(8028) := b"1111111111111111_1111111111111111_1010101000100111_0101110100000000"; -- -0.3353368639945984
	pesos_i(8029) := b"0000000000000000_0000000000000000_0011100100010001_0111111100000000"; -- 0.22292321920394897
	pesos_i(8030) := b"1111111111111111_1111111111111111_1101011010100111_0101110010000000"; -- -0.16150876879692078
	pesos_i(8031) := b"0000000000000000_0000000000000000_0000010001011100_1110001000001000"; -- 0.017042281106114388
	pesos_i(8032) := b"0000000000000000_0000000000000000_0100110111110010_1111100110000000"; -- 0.30448874831199646
	pesos_i(8033) := b"0000000000000000_0000000000000000_0001111010001110_0011101001000000"; -- 0.11935772001743317
	pesos_i(8034) := b"1111111111111111_1111111111111111_1110101111010010_0000011001000000"; -- -0.07882653176784515
	pesos_i(8035) := b"0000000000000000_0000000000000000_0000001011110101_1010110010100100"; -- 0.011561193503439426
	pesos_i(8036) := b"1111111111111111_1111111111111111_1101101101100100_1010100111000000"; -- -0.14299525320529938
	pesos_i(8037) := b"0000000000000000_0000000000000000_0000000010011011_1001100000010111"; -- 0.0023741775657981634
	pesos_i(8038) := b"1111111111111111_1111111111111111_1101011110110101_1101110010000000"; -- -0.15738126635551453
	pesos_i(8039) := b"1111111111111111_1111111111111111_1001011110000101_1100000100000000"; -- -0.40811532735824585
	pesos_i(8040) := b"0000000000000000_0000000000000000_0001110010011010_1111101100000000"; -- 0.11173981428146362
	pesos_i(8041) := b"0000000000000000_0000000000000000_0001010100011001_1100011011100000"; -- 0.0824245736002922
	pesos_i(8042) := b"0000000000000000_0000000000000000_0011011010100101_0101001100000000"; -- 0.21346014738082886
	pesos_i(8043) := b"1111111111111111_1111111111111111_1100101110001011_1001110010000000"; -- -0.20490095019340515
	pesos_i(8044) := b"1111111111111111_1111111111111111_1111001110111101_0010100100100000"; -- -0.04789488762617111
	pesos_i(8045) := b"0000000000000000_0000000000000000_0000001010001000_0100111100111000"; -- 0.0098924171179533
	pesos_i(8046) := b"1111111111111111_1111111111111111_1101110001100001_1010011000000000"; -- -0.13913500308990479
	pesos_i(8047) := b"1111111111111111_1111111111111111_1110001001010001_1000010000100000"; -- -0.11594366282224655
	pesos_i(8048) := b"1111111111111111_1111111111111111_1111111000010100_0001011100010100"; -- -0.007505948655307293
	pesos_i(8049) := b"1111111111111111_1111111111111111_1110011001111111_1010100110100000"; -- -0.09961452335119247
	pesos_i(8050) := b"1111111111111111_1111111111111111_1101011100001101_0000001000000000"; -- -0.15995776653289795
	pesos_i(8051) := b"1111111111111111_1111111111111111_1110111011101001_0100011011100000"; -- -0.06675297766923904
	pesos_i(8052) := b"1111111111111111_1111111111111111_1101101001101100_0011110011000000"; -- -0.1467859297990799
	pesos_i(8053) := b"0000000000000000_0000000000000000_0000110011111110_0111111111110000"; -- 0.05075835809111595
	pesos_i(8054) := b"0000000000000000_0000000000000000_0000001001101100_1100110001010100"; -- 0.009472628124058247
	pesos_i(8055) := b"0000000000000000_0000000000000000_0000000000101011_1110110000110001"; -- 0.0006702060345560312
	pesos_i(8056) := b"0000000000000000_0000000000000000_0001011001110001_0101110101100000"; -- 0.0876673087477684
	pesos_i(8057) := b"1111111111111111_1111111111111111_1011111110101011_0011101100000000"; -- -0.25129348039627075
	pesos_i(8058) := b"1111111111111111_1111111111111111_1101101110101001_0101100101000000"; -- -0.1419471949338913
	pesos_i(8059) := b"0000000000000000_0000000000000000_0000011110010111_0111010101101000"; -- 0.02965482510626316
	pesos_i(8060) := b"0000000000000000_0000000000000000_0010100001110110_1100111111000000"; -- 0.1580629199743271
	pesos_i(8061) := b"1111111111111111_1111111111111111_1101110011111010_1011001011000000"; -- -0.1367996484041214
	pesos_i(8062) := b"1111111111111111_1111111111111111_1110000100111101_1001001010000000"; -- -0.1201542317867279
	pesos_i(8063) := b"0000000000000000_0000000000000000_0011000101001111_0001100101000000"; -- 0.19261319935321808
	pesos_i(8064) := b"0000000000000000_0000000000000000_0001010100001010_0100001101100000"; -- 0.08218785375356674
	pesos_i(8065) := b"1111111111111111_1111111111111111_1111100101000101_0010110000010000"; -- -0.026288267225027084
	pesos_i(8066) := b"0000000000000000_0000000000000000_0000111010111011_0110101010000000"; -- 0.05754724144935608
	pesos_i(8067) := b"1111111111111111_1111111111111111_1111001001011101_0001111001110000"; -- -0.05326661840081215
	pesos_i(8068) := b"1111111111111111_1111111111111111_1111001101101111_0001011010000000"; -- -0.049086183309555054
	pesos_i(8069) := b"0000000000000000_0000000000000000_0000011111101001_0110110110110000"; -- 0.0309055857360363
	pesos_i(8070) := b"0000000000000000_0000000000000000_0000001111011001_0011110111001100"; -- 0.015033590607345104
	pesos_i(8071) := b"0000000000000000_0000000000000000_0001111110000110_1001000010000000"; -- 0.12314704060554504
	pesos_i(8072) := b"1111111111111111_1111111111111111_1100111000101000_0000110100000000"; -- -0.19470137357711792
	pesos_i(8073) := b"0000000000000000_0000000000000000_0001000101100111_1111010001000000"; -- 0.06799246370792389
	pesos_i(8074) := b"0000000000000000_0000000000000000_0001110101101010_1001111100000000"; -- 0.11490815877914429
	pesos_i(8075) := b"1111111111111111_1111111111111111_1111111011010010_0001001010111110"; -- -0.004607037175446749
	pesos_i(8076) := b"0000000000000000_0000000000000000_0001011010010110_1011110110000000"; -- 0.08823761343955994
	pesos_i(8077) := b"0000000000000000_0000000000000000_0001111001100110_1011100010100000"; -- 0.11875490099191666
	pesos_i(8078) := b"1111111111111111_1111111111111111_1110001000010100_0000000010000000"; -- -0.11688229441642761
	pesos_i(8079) := b"1111111111111111_1111111111111111_1110010101110100_1101001100000000"; -- -0.10368615388870239
	pesos_i(8080) := b"1111111111111111_1111111111111111_1111010101010000_1101000000110000"; -- -0.04173563793301582
	pesos_i(8081) := b"0000000000000000_0000000000000000_0001101001100000_1101111011000000"; -- 0.10304062068462372
	pesos_i(8082) := b"1111111111111111_1111111111111111_1111101010111111_0000010101001000"; -- -0.02052275650203228
	pesos_i(8083) := b"1111111111111111_1111111111111111_1111111001111110_1111001000001100"; -- -0.005875465460121632
	pesos_i(8084) := b"0000000000000000_0000000000000000_0001000100101000_0000011000100000"; -- 0.06701696664094925
	pesos_i(8085) := b"0000000000000000_0000000000000000_0000110010101110_1110110111100000"; -- 0.049544207751750946
	pesos_i(8086) := b"0000000000000000_0000000000000000_0001101110110110_1100010111100000"; -- 0.10825764387845993
	pesos_i(8087) := b"0000000000000000_0000000000000000_0000010001101110_0010100110100000"; -- 0.017305947840213776
	pesos_i(8088) := b"0000000000000000_0000000000000000_0000000001001111_0100011001110000"; -- 0.0012096428545191884
	pesos_i(8089) := b"0000000000000000_0000000000000000_0001010101111011_0111011111100000"; -- 0.08391522616147995
	pesos_i(8090) := b"1111111111111111_1111111111111111_1110111001011001_0010110110100000"; -- -0.06895174831151962
	pesos_i(8091) := b"1111111111111111_1111111111111111_1100111000100110_1111011101000000"; -- -0.19471792876720428
	pesos_i(8092) := b"1111111111111111_1111111111111111_1101010001010100_0000000001000000"; -- -0.1705932468175888
	pesos_i(8093) := b"1111111111111111_1111111111111111_1111100111000100_1011010001010000"; -- -0.024342279881238937
	pesos_i(8094) := b"0000000000000000_0000000000000000_0000001010011100_1110001001001000"; -- 0.010206358507275581
	pesos_i(8095) := b"1111111111111111_1111111111111111_1111010101111110_1110010000110000"; -- -0.041032541543245316
	pesos_i(8096) := b"1111111111111111_1111111111111111_1111110001010010_0110001101111100"; -- -0.014367849566042423
	pesos_i(8097) := b"0000000000000000_0000000000000000_0011000000100000_1110101010000000"; -- 0.18800225853919983
	pesos_i(8098) := b"0000000000000000_0000000000000000_0001110111011011_0010101000100000"; -- 0.11662543565034866
	pesos_i(8099) := b"1111111111111111_1111111111111111_1111001111011011_1000000000000000"; -- -0.04743194580078125
	pesos_i(8100) := b"1111111111111111_1111111111111111_1100100100001011_1111011111000000"; -- -0.2146611362695694
	pesos_i(8101) := b"0000000000000000_0000000000000000_0010011011010011_0110001010000000"; -- 0.15166297554969788
	pesos_i(8102) := b"0000000000000000_0000000000000000_0000100010010101_0110111001100000"; -- 0.033530138432979584
	pesos_i(8103) := b"0000000000000000_0000000000000000_0010100101001010_1010110011000000"; -- 0.16129569709300995
	pesos_i(8104) := b"0000000000000000_0000000000000000_0011110100111001_0110011100000000"; -- 0.23915714025497437
	pesos_i(8105) := b"1111111111111111_1111111111111111_1111000011011110_1101101010110000"; -- -0.05909951403737068
	pesos_i(8106) := b"1111111111111111_1111111111111111_1101001101010100_0111110110000000"; -- -0.1744920313358307
	pesos_i(8107) := b"0000000000000000_0000000000000000_0001010001101010_0001111001000000"; -- 0.07974423468112946
	pesos_i(8108) := b"0000000000000000_0000000000000000_0000101011000100_0011111101100000"; -- 0.04205700010061264
	pesos_i(8109) := b"1111111111111111_1111111111111111_1111110111110010_0110000011110000"; -- -0.008020345121622086
	pesos_i(8110) := b"1111111111111111_1111111111111111_1101111000111000_0011110000000000"; -- -0.13195443153381348
	pesos_i(8111) := b"1111111111111111_1111111111111111_1111101000110010_1110000000111000"; -- -0.022661196067929268
	pesos_i(8112) := b"0000000000000000_0000000000000000_0000000011000001_0000111101000111"; -- 0.0029458568897098303
	pesos_i(8113) := b"1111111111111111_1111111111111111_1101100100011101_0100001001000000"; -- -0.15189729630947113
	pesos_i(8114) := b"1111111111111111_1111111111111111_1101101001101000_0101111111000000"; -- -0.14684487879276276
	pesos_i(8115) := b"0000000000000000_0000000000000000_0001010101010010_1001100001100000"; -- 0.08329155296087265
	pesos_i(8116) := b"0000000000000000_0000000000000000_0011000010001011_0011011111000000"; -- 0.18962429463863373
	pesos_i(8117) := b"1111111111111111_1111111111111111_1110110110000101_0110001100100000"; -- -0.07218342274427414
	pesos_i(8118) := b"1111111111111111_1111111111111111_1111111110011101_1101000101100100"; -- -0.001498139463365078
	pesos_i(8119) := b"1111111111111111_1111111111111111_1111101101101101_0011110100010000"; -- -0.017864402383565903
	pesos_i(8120) := b"1111111111111111_1111111111111111_1111010110100001_1111001110010000"; -- -0.040497567504644394
	pesos_i(8121) := b"0000000000000000_0000000000000000_0010000001011110_1000000100000000"; -- 0.12644201517105103
	pesos_i(8122) := b"1111111111111111_1111111111111111_1011111010001110_1111010000000000"; -- -0.2556312084197998
	pesos_i(8123) := b"1111111111111111_1111111111111111_1110110000101001_1010011001000000"; -- -0.07748948037624359
	pesos_i(8124) := b"1111111111111111_1111111111111111_1101111010011010_1111011010000000"; -- -0.13044795393943787
	pesos_i(8125) := b"0000000000000000_0000000000000000_0010000111001000_0000110000000000"; -- 0.1319587230682373
	pesos_i(8126) := b"0000000000000000_0000000000000000_0001111111100100_0010111101000000"; -- 0.12457557022571564
	pesos_i(8127) := b"0000000000000000_0000000000000000_0000001110111001_0010011001001000"; -- 0.014543907716870308
	pesos_i(8128) := b"1111111111111111_1111111111111111_1111101101111100_1010100010111000"; -- -0.017629103735089302
	pesos_i(8129) := b"1111111111111111_1111111111111111_1111010001010000_0010011010110000"; -- -0.04565199092030525
	pesos_i(8130) := b"0000000000000000_0000000000000000_0100000110001010_1011000010000000"; -- 0.25602248311042786
	pesos_i(8131) := b"0000000000000000_0000000000000000_0101001101011010_1000011010000000"; -- 0.3256000578403473
	pesos_i(8132) := b"1111111111111111_1111111111111111_1111100100110111_1100000011000000"; -- -0.026493027806282043
	pesos_i(8133) := b"1111111111111111_1111111111111111_1011111000010011_0010100000000000"; -- -0.2575201988220215
	pesos_i(8134) := b"1111111111111111_1111111111111111_1111001001001000_0100010100010000"; -- -0.0535847507417202
	pesos_i(8135) := b"0000000000000000_0000000000000000_0001011011101101_1010000010100000"; -- 0.08956340700387955
	pesos_i(8136) := b"0000000000000000_0000000000000000_0001110011001010_0001100001100000"; -- 0.1124587282538414
	pesos_i(8137) := b"0000000000000000_0000000000000000_0010111111000010_1100001101000000"; -- 0.1865655928850174
	pesos_i(8138) := b"0000000000000000_0000000000000000_0010101100001110_1101010001000000"; -- 0.16819502413272858
	pesos_i(8139) := b"1111111111111111_1111111111111111_1101100111001011_0111110101000000"; -- -0.14923875033855438
	pesos_i(8140) := b"1111111111111111_1111111111111111_1110000000001101_0101110010000000"; -- -0.12479612231254578
	pesos_i(8141) := b"1111111111111111_1111111111111111_1111010110011100_1011000101010000"; -- -0.040577810257673264
	pesos_i(8142) := b"0000000000000000_0000000000000000_0001100100010000_1000000011000000"; -- 0.09790806472301483
	pesos_i(8143) := b"1111111111111111_1111111111111111_1100110010101010_0010010101000000"; -- -0.20052878558635712
	pesos_i(8144) := b"1111111111111111_1111111111111111_1111101100111011_1101110101101000"; -- -0.0186177846044302
	pesos_i(8145) := b"0000000000000000_0000000000000000_0001001011000000_1100110001100000"; -- 0.07325436919927597
	pesos_i(8146) := b"0000000000000000_0000000000000000_0000000011101001_1110010010110101"; -- 0.0035689298529177904
	pesos_i(8147) := b"0000000000000000_0000000000000000_0100001111111010_1001010010000000"; -- 0.26554229855537415
	pesos_i(8148) := b"1111111111111111_1111111111111111_1110110111110101_1100011101100000"; -- -0.0704684630036354
	pesos_i(8149) := b"1111111111111111_1111111111111111_1110000010000000_0100110001100000"; -- -0.12304232269525528
	pesos_i(8150) := b"0000000000000000_0000000000000000_0010000000100111_0010000101000000"; -- 0.12559707462787628
	pesos_i(8151) := b"1111111111111111_1111111111111111_1101110111010110_1000111100000000"; -- -0.13344484567642212
	pesos_i(8152) := b"0000000000000000_0000000000000000_0000000100100110_0111101011100000"; -- 0.004493407905101776
	pesos_i(8153) := b"0000000000000000_0000000000000000_0001001100110011_0110000111100000"; -- 0.07500278204679489
	pesos_i(8154) := b"1111111111111111_1111111111111111_1101001101011011_0111110001000000"; -- -0.17438529431819916
	pesos_i(8155) := b"1111111111111111_1111111111111111_1111101101001000_0100001100011000"; -- -0.0184286180883646
	pesos_i(8156) := b"1111111111111111_1111111111111111_1110001101110001_0001001000000000"; -- -0.11155593395233154
	pesos_i(8157) := b"1111111111111111_1111111111111111_1101000110010010_1001101001000000"; -- -0.1813567727804184
	pesos_i(8158) := b"1111111111111111_1111111111111111_1110011101101101_0010001101000000"; -- -0.09599094092845917
	pesos_i(8159) := b"1111111111111111_1111111111111111_1101010110000001_0101111110000000"; -- -0.16599467396736145
	pesos_i(8160) := b"0000000000000000_0000000000000000_0011010000111110_0001011010000000"; -- 0.20407238602638245
	pesos_i(8161) := b"1111111111111111_1111111111111111_1110111111101011_0101111110100000"; -- -0.06281473487615585
	pesos_i(8162) := b"0000000000000000_0000000000000000_0010000011000000_1101000011000000"; -- 0.12794212996959686
	pesos_i(8163) := b"0000000000000000_0000000000000000_0000100101100001_0000111001000000"; -- 0.03663720190525055
	pesos_i(8164) := b"1111111111111111_1111111111111111_1111010100111101_1110010010110000"; -- -0.04202433302998543
	pesos_i(8165) := b"0000000000000000_0000000000000000_0010010111011001_1110001010000000"; -- 0.14785590767860413
	pesos_i(8166) := b"1111111111111111_1111111111111111_1111001100000101_1010010001010000"; -- -0.050695162266492844
	pesos_i(8167) := b"0000000000000000_0000000000000000_0001100110010011_1001000110000000"; -- 0.09990796446800232
	pesos_i(8168) := b"0000000000000000_0000000000000000_0010110111001110_0000111110000000"; -- 0.17892548441886902
	pesos_i(8169) := b"0000000000000000_0000000000000000_0001111001000001_0001101100000000"; -- 0.11818093061447144
	pesos_i(8170) := b"0000000000000000_0000000000000000_0010001101100000_0000111011000000"; -- 0.13818447291851044
	pesos_i(8171) := b"0000000000000000_0000000000000000_0011011100101100_0110111000000000"; -- 0.2155216932296753
	pesos_i(8172) := b"0000000000000000_0000000000000000_0010001111001100_0010010001000000"; -- 0.1398337036371231
	pesos_i(8173) := b"0000000000000000_0000000000000000_0101010010110101_1101100000000000"; -- 0.330899715423584
	pesos_i(8174) := b"0000000000000000_0000000000000000_0001101101010101_0101110110000000"; -- 0.106771320104599
	pesos_i(8175) := b"1111111111111111_1111111111111111_1111001111101000_1110101001110000"; -- -0.04722723737359047
	pesos_i(8176) := b"0000000000000000_0000000000000000_0001011101111110_1100001011000000"; -- 0.09177796542644501
	pesos_i(8177) := b"0000000000000000_0000000000000000_0010010010001101_0101100000000000"; -- 0.14278173446655273
	pesos_i(8178) := b"1111111111111111_1111111111111111_1101010000101100_1100111010000000"; -- -0.17119130492210388
	pesos_i(8179) := b"1111111111111111_1111111111111111_1101110000010001_0100101000000000"; -- -0.14036118984222412
	pesos_i(8180) := b"1111111111111111_1111111111111111_1111101101010100_0001111101111000"; -- -0.018247636035084724
	pesos_i(8181) := b"1111111111111111_1111111111111111_1110101110101010_1000001110000000"; -- -0.07942941784858704
	pesos_i(8182) := b"0000000000000000_0000000000000000_0001001111010100_0011000010100000"; -- 0.0774565115571022
	pesos_i(8183) := b"1111111111111111_1111111111111111_1111111010101110_0001001111010100"; -- -0.005156288854777813
	pesos_i(8184) := b"1111111111111111_1111111111111111_1111110010101100_1111111111100100"; -- -0.012985236011445522
	pesos_i(8185) := b"1111111111111111_1111111111111111_1101010010011111_0100110100000000"; -- -0.1694442629814148
	pesos_i(8186) := b"1111111111111111_1111111111111111_1101000000100011_1110101111000000"; -- -0.1869518905878067
	pesos_i(8187) := b"0000000000000000_0000000000000000_0001011110011011_1111111110000000"; -- 0.09222409129142761
	pesos_i(8188) := b"0000000000000000_0000000000000000_0010111111010111_0100111011000000"; -- 0.18687908351421356
	pesos_i(8189) := b"1111111111111111_1111111111111111_1110000101100110_0101001100000000"; -- -0.11953240633010864
	pesos_i(8190) := b"0000000000000000_0000000000000000_0100010010011111_1100010110000000"; -- 0.26806291937828064
	pesos_i(8191) := b"0000000000000000_0000000000000000_0000000100010011_1011110101000100"; -- 0.004207448102533817
	pesos_i(8192) := b"1111111111111111_1111111111111111_0101110101110000_0111110100000000"; -- -0.6350023150444031
	pesos_i(8193) := b"1111111111111111_1111111111111111_1111111111001110_1010011000001110"; -- -0.0007530419388785958
	pesos_i(8194) := b"0000000000000000_0000000000000000_0011111101010100_0100000000000000"; -- 0.24737930297851562
	pesos_i(8195) := b"1111111111111111_1111111111111111_1111111111111101_0001011001101100"; -- -4.444000660441816e-05
	pesos_i(8196) := b"1111111111111111_1111111111111111_1101001101000111_1010100000000000"; -- -0.17468786239624023
	pesos_i(8197) := b"0000000000000000_0000000000000000_0000110000011000_0001111110100000"; -- 0.04724309593439102
	pesos_i(8198) := b"0000000000000000_0000000000000000_0000111010001111_0011111100010000"; -- 0.05687326565384865
	pesos_i(8199) := b"0000000000000000_0000000000000000_0000100010001100_1101011001010000"; -- 0.033399004489183426
	pesos_i(8200) := b"0000000000000000_0000000000000000_0010011110001001_1000000001000000"; -- 0.15444184839725494
	pesos_i(8201) := b"1111111111111111_1111111111111110_1100110100011111_1101101000000000"; -- -1.1987327337265015
	pesos_i(8202) := b"1111111111111111_1111111111111111_0110011000010101_1010111100000000"; -- -0.6012316346168518
	pesos_i(8203) := b"0000000000000000_0000000000000000_0000010000111011_1100100011101000"; -- 0.016537243500351906
	pesos_i(8204) := b"1111111111111111_1111111111111111_1111011001100100_1001111011010000"; -- -0.03752715513110161
	pesos_i(8205) := b"0000000000000000_0000000000000000_0001111101110001_0110000011100000"; -- 0.12282376736402512
	pesos_i(8206) := b"1111111111111111_1111111111111111_1010011110001101_1111110000000000"; -- -0.3454897403717041
	pesos_i(8207) := b"0000000000000000_0000000000000000_0111100001101111_0101011110000000"; -- 0.47044894099235535
	pesos_i(8208) := b"1111111111111111_1111111111111110_1111011010101000_0110000000000000"; -- -1.0364933013916016
	pesos_i(8209) := b"0000000000000000_0000000000000000_0010001011100000_1000000000000000"; -- 0.13623809814453125
	pesos_i(8210) := b"0000000000000000_0000000000000000_0000100000111100_0001010101010000"; -- 0.032166797667741776
	pesos_i(8211) := b"0000000000000000_0000000000000000_0001110101011011_0011011110100000"; -- 0.11467311531305313
	pesos_i(8212) := b"0000000000000000_0000000000000000_0111110110011100_1011010100000000"; -- 0.49067240953445435
	pesos_i(8213) := b"1111111111111111_1111111111111111_1101110010101100_1010011101000000"; -- -0.13799051940441132
	pesos_i(8214) := b"0000000000000000_0000000000000000_0111001111010101_1110010010000000"; -- 0.4524824917316437
	pesos_i(8215) := b"0000000000000000_0000000000000000_0010111011000000_1101001110000000"; -- 0.18262979388237
	pesos_i(8216) := b"1111111111111111_1111111111111111_1101111011010001_0011000101000000"; -- -0.1296204775571823
	pesos_i(8217) := b"1111111111111111_1111111111111111_1101101001101111_1010110000000000"; -- -0.14673352241516113
	pesos_i(8218) := b"1111111111111111_1111111111111111_1010100110101001_0000001010000000"; -- -0.33726486563682556
	pesos_i(8219) := b"0000000000000000_0000000000000000_0100111100000010_1001001100000000"; -- 0.308633029460907
	pesos_i(8220) := b"1111111111111111_1111111111111111_1010111010111110_1000001000000000"; -- -0.3174055814743042
	pesos_i(8221) := b"1111111111111111_1111111111111111_0010011001110100_1000011000000000"; -- -0.8497844934463501
	pesos_i(8222) := b"0000000000000000_0000000000000000_0000100010110100_1000010011110000"; -- 0.03400450572371483
	pesos_i(8223) := b"1111111111111111_1111111111111111_0110110011000110_0000010100000000"; -- -0.5751034617424011
	pesos_i(8224) := b"1111111111111111_1111111111111111_1111010100100100_1000000010010000"; -- -0.042411770671606064
	pesos_i(8225) := b"1111111111111111_1111111111111111_1001100011010101_1110000010000000"; -- -0.4029864966869354
	pesos_i(8226) := b"0000000000000000_0000000000000000_0011100100101011_0000111011000000"; -- 0.22331325709819794
	pesos_i(8227) := b"0000000000000000_0000000000000000_0011100110110010_1001100010000000"; -- 0.22538140416145325
	pesos_i(8228) := b"0000000000000000_0000000000000000_0101100101000110_1101011010000000"; -- 0.3487371504306793
	pesos_i(8229) := b"0000000000000000_0000000000000000_0010101011001001_0000001111000000"; -- 0.1671297401189804
	pesos_i(8230) := b"0000000000000000_0000000000000000_0011111011010100_1000100001000000"; -- 0.24543048441410065
	pesos_i(8231) := b"1111111111111111_1111111111111111_1110110001110010_0100111001100000"; -- -0.07638082653284073
	pesos_i(8232) := b"1111111111111111_1111111111111111_0111100000111011_0010101100000000"; -- -0.5303471684455872
	pesos_i(8233) := b"0000000000000000_0000000000000000_0100000011010011_1011000000000000"; -- 0.25323009490966797
	pesos_i(8234) := b"0000000000000000_0000000000000000_0000100101101001_1000110110000000"; -- 0.03676685690879822
	pesos_i(8235) := b"0000000000000000_0000000000000000_0111111101010010_1110000110000000"; -- 0.49735841155052185
	pesos_i(8236) := b"0000000000000000_0000000000000000_0110011110001111_1100100100000000"; -- 0.40453773736953735
	pesos_i(8237) := b"1111111111111111_1111111111111111_0110011101110100_0011000000000000"; -- -0.5958833694458008
	pesos_i(8238) := b"1111111111111111_1111111111111111_0111000111101100_1000101100000000"; -- -0.5549843907356262
	pesos_i(8239) := b"1111111111111111_1111111111111111_1110010101011010_1001011001000000"; -- -0.1040865033864975
	pesos_i(8240) := b"0000000000000000_0000000000000000_0010000101111101_1010111110000000"; -- 0.13082405924797058
	pesos_i(8241) := b"0000000000000000_0000000000000000_0000111010100011_0011100001110000"; -- 0.05717804655432701
	pesos_i(8242) := b"0000000000000000_0000000000000000_0000000010100110_0110101001101101"; -- 0.0025393024552613497
	pesos_i(8243) := b"0000000000000000_0000000000000000_0111100110000100_1111001010000000"; -- 0.47468486428260803
	pesos_i(8244) := b"0000000000000000_0000000000000000_0000110101101110_1101100010100000"; -- 0.05247262865304947
	pesos_i(8245) := b"1111111111111111_1111111111111111_1010100111100010_1111001110000000"; -- -0.3363807499408722
	pesos_i(8246) := b"1111111111111111_1111111111111111_0110001001111100_0000011100000000"; -- -0.6152949929237366
	pesos_i(8247) := b"0000000000000000_0000000000000001_0011010000011111_1111000000000000"; -- 1.2036123275756836
	pesos_i(8248) := b"1111111111111111_1111111111111111_1000110000100011_0010110100000000"; -- -0.4525882601737976
	pesos_i(8249) := b"1111111111111111_1111111111111111_1101110011001110_0001111110000000"; -- -0.13747981190681458
	pesos_i(8250) := b"1111111111111111_1111111111111111_0110010011111001_0101110100000000"; -- -0.6055700182914734
	pesos_i(8251) := b"0000000000000000_0000000000000000_0100010010110110_0010001100000000"; -- 0.26840418577194214
	pesos_i(8252) := b"0000000000000000_0000000000000000_0001001110011010_1000001001100000"; -- 0.07657637447118759
	pesos_i(8253) := b"1111111111111111_1111111111111111_1001010000111000_0000101100000000"; -- -0.42101985216140747
	pesos_i(8254) := b"0000000000000000_0000000000000000_0001101100010110_0100001001000000"; -- 0.10580839216709137
	pesos_i(8255) := b"0000000000000000_0000000000000000_0100001110001010_0101101100000000"; -- 0.26382988691329956
	pesos_i(8256) := b"1111111111111111_1111111111111111_1110001100010011_0110011111100000"; -- -0.11298514157533646
	pesos_i(8257) := b"0000000000000000_0000000000000000_0001011110101111_1011000101100000"; -- 0.09252461045980453
	pesos_i(8258) := b"0000000000000000_0000000000000000_0001001011101010_1110010110000000"; -- 0.07389673590660095
	pesos_i(8259) := b"1111111111111111_1111111111111111_0011101111100011_0110101100000000"; -- -0.7660611271858215
	pesos_i(8260) := b"1111111111111111_1111111111111111_1110110010100010_1001001101000000"; -- -0.07564429938793182
	pesos_i(8261) := b"1111111111111111_1111111111111111_1011011101101110_0001000100000000"; -- -0.2834767699241638
	pesos_i(8262) := b"0000000000000000_0000000000000000_0011100001010100_1110101111000000"; -- 0.2200457900762558
	pesos_i(8263) := b"0000000000000000_0000000000000000_0101011111010111_0111111010000000"; -- 0.3431319296360016
	pesos_i(8264) := b"1111111111111111_1111111111111111_1010011001001011_1010101000000000"; -- -0.3504079580307007
	pesos_i(8265) := b"1111111111111111_1111111111111111_1111001010011000_1100110010010000"; -- -0.052355971187353134
	pesos_i(8266) := b"1111111111111111_1111111111111111_1110111111000000_0001001001000000"; -- -0.06347547471523285
	pesos_i(8267) := b"1111111111111111_1111111111111111_1111111100101100_1001011101001010"; -- -0.0032258457504212856
	pesos_i(8268) := b"0000000000000000_0000000000000000_0001111011101001_1011100100100000"; -- 0.12075383216142654
	pesos_i(8269) := b"0000000000000000_0000000000000000_0101001110111001_0111010000000000"; -- 0.32704854011535645
	pesos_i(8270) := b"1111111111111111_1111111111111111_0010101101010000_0001001100000000"; -- -0.8308094143867493
	pesos_i(8271) := b"1111111111111111_1111111111111111_1100100100111100_1001000010000000"; -- -0.21391960978507996
	pesos_i(8272) := b"1111111111111111_1111111111111111_1000011000011101_0111101100000000"; -- -0.4761126637458801
	pesos_i(8273) := b"0000000000000000_0000000000000000_0111100010000100_0000011010000000"; -- 0.47076454758644104
	pesos_i(8274) := b"1111111111111111_1111111111111111_1111000001011010_0001000011010000"; -- -0.061125706881284714
	pesos_i(8275) := b"1111111111111111_1111111111111111_1101001000100011_0101111001000000"; -- -0.17914782464504242
	pesos_i(8276) := b"0000000000000000_0000000000000000_0110110100011100_1110000100000000"; -- 0.42622190713882446
	pesos_i(8277) := b"1111111111111111_1111111111111111_0111010111101100_1100011000000000"; -- -0.5393558740615845
	pesos_i(8278) := b"1111111111111111_1111111111111111_0101110111111011_1000110000000000"; -- -0.632880449295044
	pesos_i(8279) := b"0000000000000000_0000000000000000_0100011011011110_1111001110000000"; -- 0.2768394649028778
	pesos_i(8280) := b"0000000000000000_0000000000000000_0001001110100010_0010011111000000"; -- 0.07669304311275482
	pesos_i(8281) := b"0000000000000000_0000000000000000_0000010110001110_0000101001100000"; -- 0.021698616445064545
	pesos_i(8282) := b"0000000000000000_0000000000000000_0010011010110101_1110111111000000"; -- 0.1512136310338974
	pesos_i(8283) := b"1111111111111111_1111111111111111_1111110101010110_1000010111011000"; -- -0.010398516431450844
	pesos_i(8284) := b"0000000000000000_0000000000000000_0000011101100001_1110000000111000"; -- 0.028837217018008232
	pesos_i(8285) := b"1111111111111111_1111111111111111_1011111100010100_0000000110000000"; -- -0.25360098481178284
	pesos_i(8286) := b"1111111111111111_1111111111111111_1101010100110110_0101100000000000"; -- -0.16713953018188477
	pesos_i(8287) := b"0000000000000000_0000000000000000_0101000001111100_1011000010000000"; -- 0.31440261006355286
	pesos_i(8288) := b"1111111111111111_1111111111111111_1011110011111010_1111100010000000"; -- -0.2617954909801483
	pesos_i(8289) := b"1111111111111111_1111111111111111_1001001110111000_1001100100000000"; -- -0.42296451330184937
	pesos_i(8290) := b"0000000000000000_0000000000000000_0110011001000111_0100011100000000"; -- 0.39952510595321655
	pesos_i(8291) := b"1111111111111111_1111111111111111_1110011000001111_1001000100100000"; -- -0.10132496803998947
	pesos_i(8292) := b"1111111111111111_1111111111111111_1011001001001010_0010001110000000"; -- -0.3035562336444855
	pesos_i(8293) := b"1111111111111111_1111111111111111_0111100111000101_0000100000000000"; -- -0.5243372917175293
	pesos_i(8294) := b"1111111111111111_1111111111111111_0111101110111000_1010011000000000"; -- -0.5167137384414673
	pesos_i(8295) := b"0000000000000000_0000000000000000_0110001011000111_1100001100000000"; -- 0.3858606219291687
	pesos_i(8296) := b"0000000000000000_0000000000000000_0010010110111111_1101100000000000"; -- 0.14745855331420898
	pesos_i(8297) := b"0000000000000000_0000000000000000_0010100111100011_0110000000000000"; -- 0.16362571716308594
	pesos_i(8298) := b"1111111111111111_1111111111111111_1010011101101011_1000100100000000"; -- -0.34601539373397827
	pesos_i(8299) := b"0000000000000000_0000000000000000_0010101001000100_1110001101000000"; -- 0.1651136428117752
	pesos_i(8300) := b"1111111111111111_1111111111111111_1110101011110001_0000000010000000"; -- -0.08226010203361511
	pesos_i(8301) := b"1111111111111111_1111111111111111_1101111010011011_1111110110000000"; -- -0.13043227791786194
	pesos_i(8302) := b"1111111111111111_1111111111111111_1011110001110010_0110100010000000"; -- -0.26387926936149597
	pesos_i(8303) := b"0000000000000000_0000000000000000_0011011001111000_0110100001000000"; -- 0.21277476847171783
	pesos_i(8304) := b"1111111111111111_1111111111111111_1110101110011000_0011000001100000"; -- -0.07970903068780899
	pesos_i(8305) := b"0000000000000000_0000000000000000_0110101100110111_0110111100000000"; -- 0.41881459951400757
	pesos_i(8306) := b"1111111111111111_1111111111111111_0100010111010011_0101111100000000"; -- -0.7272434830665588
	pesos_i(8307) := b"1111111111111111_1111111111111111_0111100101010000_1011111000000000"; -- -0.5261117219924927
	pesos_i(8308) := b"0000000000000000_0000000000000000_0001100110110011_1100110010000000"; -- 0.10039976239204407
	pesos_i(8309) := b"0000000000000000_0000000000000000_0110010101101001_1110011010000000"; -- 0.3961471617221832
	pesos_i(8310) := b"1111111111111111_1111111111111111_1111000000111100_0011110110100000"; -- -0.06158079952001572
	pesos_i(8311) := b"0000000000000000_0000000000000000_0010101001010011_0100000011000000"; -- 0.1653328388929367
	pesos_i(8312) := b"0000000000000000_0000000000000000_0011011111010000_0110010110000000"; -- 0.2180236279964447
	pesos_i(8313) := b"0000000000000000_0000000000000000_0000100010100000_1100100100010000"; -- 0.03370339050889015
	pesos_i(8314) := b"1111111111111111_1111111111111111_0110010111100011_1111010100000000"; -- -0.6019904017448425
	pesos_i(8315) := b"1111111111111111_1111111111111111_1010011000001100_0110000110000000"; -- -0.3513735830783844
	pesos_i(8316) := b"0000000000000000_0000000000000000_0000000011001010_1111100001100110"; -- 0.0030970810912549496
	pesos_i(8317) := b"1111111111111111_1111111111111111_1110111101000110_1100001000000000"; -- -0.06532657146453857
	pesos_i(8318) := b"0000000000000000_0000000000000000_0011101100100101_1111100110000000"; -- 0.23104819655418396
	pesos_i(8319) := b"1111111111111111_1111111111111111_1111110111011101_0101010010011000"; -- -0.008341515436768532
	pesos_i(8320) := b"1111111111111111_1111111111111111_1111101110111100_0110100100001000"; -- -0.016656337305903435
	pesos_i(8321) := b"0000000000000000_0000000000000000_0000001111010110_1111101000111100"; -- 0.014999045990407467
	pesos_i(8322) := b"0000000000000000_0000000000000000_0110010100100100_0001101000000000"; -- 0.39508211612701416
	pesos_i(8323) := b"1111111111111111_1111111111111111_1100001000110100_1100111100000000"; -- -0.2413817048072815
	pesos_i(8324) := b"0000000000000000_0000000000000000_0000101011111001_0011110111000000"; -- 0.04286561906337738
	pesos_i(8325) := b"1111111111111111_1111111111111111_1101110001001100_0101110110000000"; -- -0.1394597589969635
	pesos_i(8326) := b"0000000000000000_0000000000000000_0111000000111011_1010101100000000"; -- 0.4384104609489441
	pesos_i(8327) := b"1111111111111111_1111111111111111_1110001111010111_1011001001000000"; -- -0.10998998582363129
	pesos_i(8328) := b"0000000000000000_0000000000000000_0110000010100010_1001011010000000"; -- 0.3774808943271637
	pesos_i(8329) := b"1111111111111111_1111111111111111_1001111101001001_0000110010000000"; -- -0.3777916133403778
	pesos_i(8330) := b"1111111111111111_1111111111111111_0110100001011000_0111100000000000"; -- -0.592400074005127
	pesos_i(8331) := b"1111111111111111_1111111111111111_1010101000000001_1011010100000000"; -- -0.33591145277023315
	pesos_i(8332) := b"0000000000000000_0000000000000000_0101010100001010_0011100100000000"; -- 0.3321872353553772
	pesos_i(8333) := b"1111111111111111_1111111111111111_1110000001110000_0100101010000000"; -- -0.12328657507896423
	pesos_i(8334) := b"0000000000000000_0000000000000000_0110111000100110_1111100100000000"; -- 0.4302821755409241
	pesos_i(8335) := b"0000000000000000_0000000000000000_0010011111010111_0000111111000000"; -- 0.1556253284215927
	pesos_i(8336) := b"0000000000000000_0000000000000000_0011110010001110_0111000110000000"; -- 0.236548513174057
	pesos_i(8337) := b"1111111111111111_1111111111111111_0111111110000011_1011010000000000"; -- -0.5018966197967529
	pesos_i(8338) := b"0000000000000000_0000000000000000_0100110110000011_1100111000000000"; -- 0.30279242992401123
	pesos_i(8339) := b"1111111111111111_1111111111111111_1001000100110001_1111011010000000"; -- -0.43283137679100037
	pesos_i(8340) := b"1111111111111111_1111111111111111_0111100100100110_1011000000000000"; -- -0.5267534255981445
	pesos_i(8341) := b"1111111111111111_1111111111111111_1011101100101101_1010101100000000"; -- -0.2688344120979309
	pesos_i(8342) := b"0000000000000000_0000000000000000_0100010000001011_0100010100000000"; -- 0.265796959400177
	pesos_i(8343) := b"1111111111111111_1111111111111111_1101101100100110_1101111011000000"; -- -0.14393813908100128
	pesos_i(8344) := b"1111111111111111_1111111111111111_1000001110010000_1001000010000000"; -- -0.48607537150382996
	pesos_i(8345) := b"0000000000000000_0000000000000000_0100010010100001_0110001110000000"; -- 0.26808759570121765
	pesos_i(8346) := b"0000000000000000_0000000000000000_0000101110100101_0010010011100000"; -- 0.04548864811658859
	pesos_i(8347) := b"1111111111111111_1111111111111111_1100110110111001_1000011011000000"; -- -0.19638784229755402
	pesos_i(8348) := b"1111111111111111_1111111111111111_1000111110000100_1101001000000000"; -- -0.43937957286834717
	pesos_i(8349) := b"0000000000000000_0000000000000000_0011000110000001_0100010110000000"; -- 0.1933787763118744
	pesos_i(8350) := b"1111111111111111_1111111111111111_1010001010000101_1111110100000000"; -- -0.3651430010795593
	pesos_i(8351) := b"0000000000000000_0000000000000000_0000100101111010_1111111110010000"; -- 0.03703305497765541
	pesos_i(8352) := b"1111111111111111_1111111111111111_0100100010000111_0101011100000000"; -- -0.716684877872467
	pesos_i(8353) := b"1111111111111111_1111111111111111_1110111000111001_0110011100100000"; -- -0.06943660229444504
	pesos_i(8354) := b"0000000000000000_0000000000000000_0000001111010110_0000110100010100"; -- 0.014984910376369953
	pesos_i(8355) := b"1111111111111111_1111111111111111_1011010001110101_0001000000000000"; -- -0.2950887680053711
	pesos_i(8356) := b"0000000000000000_0000000000000000_0010111000100101_0110101001000000"; -- 0.18025840818881989
	pesos_i(8357) := b"0000000000000000_0000000000000000_0000111101101101_0001111110100000"; -- 0.06025884300470352
	pesos_i(8358) := b"0000000000000000_0000000000000000_0000111000110110_0100101011000000"; -- 0.05551593005657196
	pesos_i(8359) := b"1111111111111111_1111111111111111_1100110001100110_0000100001000000"; -- -0.2015681117773056
	pesos_i(8360) := b"1111111111111111_1111111111111111_1110111110000110_0111101101100000"; -- -0.06435421854257584
	pesos_i(8361) := b"0000000000000000_0000000000000000_0101011000100101_0010100110000000"; -- 0.3365045487880707
	pesos_i(8362) := b"1111111111111111_1111111111111111_1110100100011011_0000000110100000"; -- -0.08943166583776474
	pesos_i(8363) := b"1111111111111111_1111111111111111_1111101100100011_1011101000100000"; -- -0.01898609846830368
	pesos_i(8364) := b"0000000000000000_0000000000000000_0011001110101010_0110101100000000"; -- 0.20181912183761597
	pesos_i(8365) := b"0000000000000000_0000000000000000_0010110000111111_1100111100000000"; -- 0.172848641872406
	pesos_i(8366) := b"1111111111111111_1111111111111111_1101011011100011_0110011111000000"; -- -0.16059257090091705
	pesos_i(8367) := b"1111111111111111_1111111111111111_1111011100111100_0000010110100000"; -- -0.03424038738012314
	pesos_i(8368) := b"0000000000000000_0000000000000000_0011111010011000_1010100001000000"; -- 0.24451686441898346
	pesos_i(8369) := b"1111111111111111_1111111111111111_0100010111100001_1111011100000000"; -- -0.727020800113678
	pesos_i(8370) := b"0000000000000000_0000000000000000_0011010001101010_1101100010000000"; -- 0.20475533604621887
	pesos_i(8371) := b"1111111111111111_1111111111111111_1011010110010100_1111000010000000"; -- -0.2906961143016815
	pesos_i(8372) := b"0000000000000000_0000000000000000_0001100100010011_0110100111000000"; -- 0.0979524701833725
	pesos_i(8373) := b"0000000000000000_0000000000000000_0101001000011000_1000100010000000"; -- 0.32068684697151184
	pesos_i(8374) := b"0000000000000000_0000000000000000_0101011110111110_1000001000000000"; -- 0.3427506685256958
	pesos_i(8375) := b"1111111111111111_1111111111111111_1100010001110011_0101010111000000"; -- -0.232615128159523
	pesos_i(8376) := b"1111111111111111_1111111111111111_0110001010101011_0011011000000000"; -- -0.6145750284194946
	pesos_i(8377) := b"1111111111111111_1111111111111111_1100010100000000_0001110000000000"; -- -0.2304670810699463
	pesos_i(8378) := b"1111111111111111_1111111111111111_1010110011010001_1000101010000000"; -- -0.3249276578426361
	pesos_i(8379) := b"1111111111111111_1111111111111111_0101101101111000_1101010000000000"; -- -0.6426875591278076
	pesos_i(8380) := b"0000000000000000_0000000000000000_0011011001001111_0010010111000000"; -- 0.21214519441127777
	pesos_i(8381) := b"0000000000000000_0000000000000000_0001101001011110_1111110101000000"; -- 0.10301192104816437
	pesos_i(8382) := b"0000000000000000_0000000000000000_0011100101101001_0101100010000000"; -- 0.22426369786262512
	pesos_i(8383) := b"0000000000000000_0000000000000000_0111100000100010_1010110110000000"; -- 0.46927914023399353
	pesos_i(8384) := b"0000000000000000_0000000000000000_0101101011001001_0001011100000000"; -- 0.35463088750839233
	pesos_i(8385) := b"1111111111111111_1111111111111111_1010111100111101_0001100010000000"; -- -0.3154740035533905
	pesos_i(8386) := b"1111111111111111_1111111111111111_1100001010000011_0111001000000000"; -- -0.2401818037033081
	pesos_i(8387) := b"1111111111111111_1111111111111111_1000001000001011_0001010010000000"; -- -0.4920184314250946
	pesos_i(8388) := b"0000000000000000_0000000000000000_0011000101110100_1000010000000000"; -- 0.19318413734436035
	pesos_i(8389) := b"1111111111111111_1111111111111111_1101111010110101_1100101000000000"; -- -0.13003861904144287
	pesos_i(8390) := b"1111111111111111_1111111111111111_1110101011010000_1011101111100000"; -- -0.08275247365236282
	pesos_i(8391) := b"1111111111111111_1111111111111111_1110111011001111_1010000011100000"; -- -0.06714434176683426
	pesos_i(8392) := b"0000000000000000_0000000000000000_0000011010001110_1010010100001000"; -- 0.02561408467590809
	pesos_i(8393) := b"1111111111111111_1111111111111111_0110011001110000_1000000100000000"; -- -0.599845826625824
	pesos_i(8394) := b"0000000000000000_0000000000000000_0010110011101101_1101010011000000"; -- 0.17550401389598846
	pesos_i(8395) := b"1111111111111111_1111111111111111_1111111110110000_1101000011000100"; -- -0.0012082598404958844
	pesos_i(8396) := b"0000000000000000_0000000000000000_0000010111101101_0110100111111000"; -- 0.023153899237513542
	pesos_i(8397) := b"0000000000000000_0000000000000000_0001011111110011_0101011001100000"; -- 0.09355678409337997
	pesos_i(8398) := b"0000000000000000_0000000000000000_0110000101000100_1000001100000000"; -- 0.3799516558647156
	pesos_i(8399) := b"1111111111111111_1111111111111111_1001101110010010_0001101110000000"; -- -0.3923018276691437
	pesos_i(8400) := b"0000000000000000_0000000000000000_0011111001101111_0101100101000000"; -- 0.2438865453004837
	pesos_i(8401) := b"1111111111111111_1111111111111111_1110100000010100_0111000111000000"; -- -0.0934380441904068
	pesos_i(8402) := b"1111111111111111_1111111111111111_1000000000011100_0001110000000000"; -- -0.4995710849761963
	pesos_i(8403) := b"0000000000000000_0000000000000000_0011010011010111_1111100011000000"; -- 0.20642046630382538
	pesos_i(8404) := b"0000000000000000_0000000000000000_0010000011001100_0010110011000000"; -- 0.1281154602766037
	pesos_i(8405) := b"0000000000000000_0000000000000000_0001111111111010_1100100110100000"; -- 0.12492046505212784
	pesos_i(8406) := b"0000000000000000_0000000000000000_0100000011001010_1101001100000000"; -- 0.2530948519706726
	pesos_i(8407) := b"1111111111111111_1111111111111111_0110100110011010_1101100000000000"; -- -0.5874810218811035
	pesos_i(8408) := b"1111111111111111_1111111111111111_1101100001110010_0000100011000000"; -- -0.15450997650623322
	pesos_i(8409) := b"1111111111111111_1111111111111111_1110100011100011_1000101001100000"; -- -0.0902780070900917
	pesos_i(8410) := b"1111111111111111_1111111111111111_1110001110010110_0111100011000000"; -- -0.11098523437976837
	pesos_i(8411) := b"0000000000000000_0000000000000000_0011100011010110_1100001001000000"; -- 0.22202695906162262
	pesos_i(8412) := b"0000000000000000_0000000000000000_1000010111110111_0011101000000000"; -- 0.5233036279678345
	pesos_i(8413) := b"0000000000000000_0000000000000000_0010101100011100_0100100011000000"; -- 0.1684003323316574
	pesos_i(8414) := b"1111111111111111_1111111111111111_1010111100011010_0100101010000000"; -- -0.31600508093833923
	pesos_i(8415) := b"0000000000000000_0000000000000000_0011100000110100_0011100000000000"; -- 0.21954679489135742
	pesos_i(8416) := b"1111111111111111_1111111111111111_0001011111110001_0110011100000000"; -- -0.9064727425575256
	pesos_i(8417) := b"0000000000000000_0000000000000000_0110011100100000_1001001000000000"; -- 0.4028407335281372
	pesos_i(8418) := b"1111111111111111_1111111111111111_0111001101001011_1110001100000000"; -- -0.5496233105659485
	pesos_i(8419) := b"0000000000000000_0000000000000000_0101010010000100_0010010010000000"; -- 0.3301413357257843
	pesos_i(8420) := b"1111111111111111_1111111111111111_0011001001001011_1010010000000000"; -- -0.8035333156585693
	pesos_i(8421) := b"1111111111111111_1111111111111111_0110111001010000_0001110100000000"; -- -0.5690900683403015
	pesos_i(8422) := b"1111111111111111_1111111111111111_0111100001100001_1100011000000000"; -- -0.529758095741272
	pesos_i(8423) := b"0000000000000000_0000000000000000_0000100011011011_0100011101110000"; -- 0.03459593281149864
	pesos_i(8424) := b"1111111111111111_1111111111111111_1011001010110010_1100001110000000"; -- -0.3019597828388214
	pesos_i(8425) := b"1111111111111111_1111111111111111_1111110011001100_1010001101000000"; -- -0.012502476572990417
	pesos_i(8426) := b"0000000000000000_0000000000000000_0011100000000100_1110100000000000"; -- 0.2188248634338379
	pesos_i(8427) := b"1111111111111111_1111111111111111_1100000100001100_1001001010000000"; -- -0.2459019124507904
	pesos_i(8428) := b"1111111111111111_1111111111111111_1111001111100000_1110001011000000"; -- -0.04734976589679718
	pesos_i(8429) := b"1111111111111111_1111111111111111_1110011101101001_1010101010000000"; -- -0.0960439145565033
	pesos_i(8430) := b"0000000000000000_0000000000000000_0000010110111100_1111100101010000"; -- 0.022414762526750565
	pesos_i(8431) := b"0000000000000000_0000000000000000_0101100101011001_1001100000000000"; -- 0.34902334213256836
	pesos_i(8432) := b"1111111111111111_1111111111111111_1101110101001010_1010001100000000"; -- -0.1355798840522766
	pesos_i(8433) := b"1111111111111111_1111111111111111_1100111011110001_0001011000000000"; -- -0.19163382053375244
	pesos_i(8434) := b"0000000000000000_0000000000000000_1001110100001100_0001101100000000"; -- 0.6134659647941589
	pesos_i(8435) := b"1111111111111111_1111111111111111_1000110000110110_1101101000000000"; -- -0.45228803157806396
	pesos_i(8436) := b"0000000000000000_0000000000000000_1000100011011100_0101100000000000"; -- 0.5346121788024902
	pesos_i(8437) := b"0000000000000000_0000000000000000_1000010100011010_1011010000000000"; -- 0.5199387073516846
	pesos_i(8438) := b"1111111111111111_1111111111111111_0000110110100001_1111110000000000"; -- -0.9467470645904541
	pesos_i(8439) := b"0000000000000000_0000000000000000_0000010000100011_1000010110011000"; -- 0.016167020425200462
	pesos_i(8440) := b"1111111111111111_1111111111111111_0101010100100011_0111101100000000"; -- -0.6674273610115051
	pesos_i(8441) := b"1111111111111111_1111111111111111_1111010100100010_1010100110010000"; -- -0.04243984445929527
	pesos_i(8442) := b"0000000000000000_0000000000000000_0010001010111110_0010110100000000"; -- 0.1357143521308899
	pesos_i(8443) := b"1111111111111111_1111111111111111_1000001110011111_1111010010000000"; -- -0.4858405292034149
	pesos_i(8444) := b"1111111111111111_1111111111111111_1000010111110000_0000010100000000"; -- -0.4768063426017761
	pesos_i(8445) := b"1111111111111111_1111111111111111_1100111100011100_0111011001000000"; -- -0.1909719556570053
	pesos_i(8446) := b"0000000000000000_0000000000000000_0101000110101100_1011111100000000"; -- 0.3190421462059021
	pesos_i(8447) := b"1111111111111111_1111111111111111_1111100110000001_0111000000111000"; -- -0.02536867745220661
	pesos_i(8448) := b"1111111111111111_1111111111111111_1100111111111011_1010100010000000"; -- -0.18756625056266785
	pesos_i(8449) := b"0000000000000000_0000000000000000_0100101100010001_1010000010000000"; -- 0.29323771595954895
	pesos_i(8450) := b"0000000000000000_0000000000000000_0001111111110010_0111011100100000"; -- 0.12479347735643387
	pesos_i(8451) := b"0000000000000000_0000000000000000_0011000100011101_1011000010000000"; -- 0.19185927510261536
	pesos_i(8452) := b"1111111111111111_1111111111111111_1100101011111111_1101011100000000"; -- -0.2070336937904358
	pesos_i(8453) := b"0000000000000000_0000000000000000_0110011101110100_1001110100000000"; -- 0.40412312746047974
	pesos_i(8454) := b"0000000000000000_0000000000000000_0010111110110110_0011100000000000"; -- 0.18637418746948242
	pesos_i(8455) := b"0000000000000000_0000000000000000_0110101011111011_0000101110000000"; -- 0.4178931415081024
	pesos_i(8456) := b"0000000000000000_0000000000000000_0000010011011010_1111011110101000"; -- 0.018966177478432655
	pesos_i(8457) := b"0000000000000000_0000000000000000_0000100111110110_0110111011100000"; -- 0.03891652077436447
	pesos_i(8458) := b"1111111111111111_1111111111111111_0111010000010110_0001010100000000"; -- -0.5465380549430847
	pesos_i(8459) := b"1111111111111111_1111111111111111_1010001110011110_0111100010000000"; -- -0.36086317896842957
	pesos_i(8460) := b"1111111111111111_1111111111111111_1111111100101101_0100001110111110"; -- -0.0032155667431652546
	pesos_i(8461) := b"1111111111111111_1111111111111111_1111001000000000_0101110110110000"; -- -0.054681915789842606
	pesos_i(8462) := b"1111111111111111_1111111111111111_1110001010010010_0011100100000000"; -- -0.1149563193321228
	pesos_i(8463) := b"0000000000000000_0000000000000000_0110100101000010_1110001000000000"; -- 0.41117680072784424
	pesos_i(8464) := b"1111111111111111_1111111111111111_1100111101011001_1100001111000000"; -- -0.19003655016422272
	pesos_i(8465) := b"0000000000000000_0000000000000000_0000000010101110_1001101110000101"; -- 0.0026642989832907915
	pesos_i(8466) := b"1111111111111111_1111111111111111_1011001001000001_1001001100000000"; -- -0.3036869168281555
	pesos_i(8467) := b"1111111111111111_1111111111111111_0011011000101011_1011010000000000"; -- -0.7883956432342529
	pesos_i(8468) := b"0000000000000000_0000000000000000_0000001100110010_1100010111001000"; -- 0.012493478134274483
	pesos_i(8469) := b"0000000000000000_0000000000000000_0101101011110100_1001010110000000"; -- 0.3552945554256439
	pesos_i(8470) := b"0000000000000000_0000000000000000_0100111000001111_0110110000000000"; -- 0.30492281913757324
	pesos_i(8471) := b"1111111111111111_1111111111111111_1101000010101001_0110100000000000"; -- -0.18491506576538086
	pesos_i(8472) := b"0000000000000000_0000000000000000_0000101110011000_1000101110100000"; -- 0.045296408236026764
	pesos_i(8473) := b"1111111111111111_1111111111111111_0101110010110111_1100001000000000"; -- -0.6378210783004761
	pesos_i(8474) := b"0000000000000000_0000000000000000_0010100000001000_0110000001000000"; -- 0.15637780725955963
	pesos_i(8475) := b"1111111111111111_1111111111111111_1000000110100001_1000111000000000"; -- -0.4936286211013794
	pesos_i(8476) := b"1111111111111111_1111111111111111_0111111011011011_1011110000000000"; -- -0.5044596195220947
	pesos_i(8477) := b"0000000000000000_0000000000000000_0110100111000011_1001010010000000"; -- 0.41314056515693665
	pesos_i(8478) := b"0000000000000000_0000000000000000_0100110011100001_0010001010000000"; -- 0.30031028389930725
	pesos_i(8479) := b"0000000000000000_0000000000000001_0000101010011011_1010111000000000"; -- 1.0414379835128784
	pesos_i(8480) := b"1111111111111111_1111111111111111_0100101110010001_1000001000000000"; -- -0.7048109769821167
	pesos_i(8481) := b"1111111111111111_1111111111111111_0010111100001010_1001110100000000"; -- -0.8162443041801453
	pesos_i(8482) := b"0000000000000000_0000000000000000_0110100010101010_0010111010000000"; -- 0.40884676575660706
	pesos_i(8483) := b"1111111111111111_1111111111111111_0110001101000010_0101110100000000"; -- -0.6122686266899109
	pesos_i(8484) := b"0000000000000000_0000000000000000_0001000110011111_1010100101000000"; -- 0.06884248554706573
	pesos_i(8485) := b"1111111111111111_1111111111111111_1010110010011111_1110001010000000"; -- -0.3256853520870209
	pesos_i(8486) := b"1111111111111111_1111111111111111_1101110110011100_1110001100000000"; -- -0.134324848651886
	pesos_i(8487) := b"0000000000000000_0000000000000000_0010110101100100_1110101000000000"; -- 0.17732107639312744
	pesos_i(8488) := b"0000000000000000_0000000000000000_0011111111101111_0101111001000000"; -- 0.24974621832370758
	pesos_i(8489) := b"1111111111111111_1111111111111111_1101111101001101_0011110000000000"; -- -0.12772774696350098
	pesos_i(8490) := b"0000000000000000_0000000000000000_0101011110011110_1110010000000000"; -- 0.3422682285308838
	pesos_i(8491) := b"1111111111111111_1111111111111111_1110100100100110_1001100110100000"; -- -0.08925475925207138
	pesos_i(8492) := b"1111111111111111_1111111111111111_1100100000001101_1101010110000000"; -- -0.21853891015052795
	pesos_i(8493) := b"1111111111111111_1111111111111111_1110011001111010_1100101010000000"; -- -0.09968885779380798
	pesos_i(8494) := b"1111111111111111_1111111111111111_1100101100111000_1100111010000000"; -- -0.20616444945335388
	pesos_i(8495) := b"0000000000000000_0000000000000000_0001000101110110_0111000101000000"; -- 0.06821353733539581
	pesos_i(8496) := b"1111111111111111_1111111111111111_1001101111111111_0101100010000000"; -- -0.3906349837779999
	pesos_i(8497) := b"1111111111111111_1111111111111111_1101100110100101_0100000011000000"; -- -0.1498221904039383
	pesos_i(8498) := b"1111111111111111_1111111111111110_1111101000011100_0010100000000000"; -- -1.023007869720459
	pesos_i(8499) := b"0000000000000000_0000000000000000_0001110001011000_1101000100000000"; -- 0.11073023080825806
	pesos_i(8500) := b"0000000000000000_0000000000000000_0000101110110010_1011101101010000"; -- 0.04569597914814949
	pesos_i(8501) := b"1111111111111111_1111111111111111_1101010001011001_1001111110000000"; -- -0.17050746083259583
	pesos_i(8502) := b"0000000000000000_0000000000000000_0000010000110010_1000111110011000"; -- 0.016396498307585716
	pesos_i(8503) := b"1111111111111111_1111111111111111_1000000100100001_1110010100000000"; -- -0.49557656049728394
	pesos_i(8504) := b"1111111111111111_1111111111111111_1001100111010010_0110101010000000"; -- -0.3991330564022064
	pesos_i(8505) := b"1111111111111111_1111111111111111_1001010111011101_0011000010000000"; -- -0.4145936667919159
	pesos_i(8506) := b"1111111111111111_1111111111111111_1001101010001110_1101101000000000"; -- -0.39625775814056396
	pesos_i(8507) := b"1111111111111111_1111111111111111_1011100010111101_0110000000000000"; -- -0.27836036682128906
	pesos_i(8508) := b"0000000000000000_0000000000000000_0001001000100001_0111000000000000"; -- 0.07082271575927734
	pesos_i(8509) := b"0000000000000000_0000000000000000_0101001000001110_1101111100000000"; -- 0.3205394148826599
	pesos_i(8510) := b"0000000000000000_0000000000000000_0100111001001000_1010011010000000"; -- 0.3057960569858551
	pesos_i(8511) := b"0000000000000000_0000000000000000_0011101000010101_0100000101000000"; -- 0.2268868237733841
	pesos_i(8512) := b"1111111111111111_1111111111111111_1010000111011100_1110000000000000"; -- -0.3677234649658203
	pesos_i(8513) := b"0000000000000000_0000000000000000_1101110100001110_0101001000000000"; -- 0.8634997606277466
	pesos_i(8514) := b"0000000000000000_0000000000000000_0000101011010001_0000011001100000"; -- 0.04225196689367294
	pesos_i(8515) := b"1111111111111111_1111111111111111_1010010000100000_0011000110000000"; -- -0.3588837683200836
	pesos_i(8516) := b"0000000000000000_0000000000000000_0101000011001101_0011100110000000"; -- 0.3156314790248871
	pesos_i(8517) := b"0000000000000000_0000000000000000_0001101101110000_0110011000100000"; -- 0.10718382149934769
	pesos_i(8518) := b"0000000000000000_0000000000000000_0111110010101110_0110001000000000"; -- 0.487035870552063
	pesos_i(8519) := b"0000000000000000_0000000000000000_0101100101111000_0000110010000000"; -- 0.3494880497455597
	pesos_i(8520) := b"1111111111111111_1111111111111111_0000011101011111_1001011100000000"; -- -0.9711976647377014
	pesos_i(8521) := b"1111111111111111_1111111111111110_0111010100101011_0011100000000000"; -- -1.542309284210205
	pesos_i(8522) := b"0000000000000000_0000000000000000_0101000110010010_0011100000000000"; -- 0.3186373710632324
	pesos_i(8523) := b"1111111111111111_1111111111111111_1110000011101011_0001110000000000"; -- -0.12141251564025879
	pesos_i(8524) := b"0000000000000000_0000000000000000_0100000110111001_0011100010000000"; -- 0.2567324936389923
	pesos_i(8525) := b"1111111111111111_1111111111111111_1110000100100110_1110101010100000"; -- -0.12049993127584457
	pesos_i(8526) := b"0000000000000000_0000000000000000_0111111110111010_0110110010000000"; -- 0.49893835186958313
	pesos_i(8527) := b"0000000000000000_0000000000000000_0101010101100101_0010111000000000"; -- 0.33357512950897217
	pesos_i(8528) := b"1111111111111111_1111111111111111_1110011011010110_0010010010000000"; -- -0.0982949435710907
	pesos_i(8529) := b"1111111111111111_1111111111111111_1001111011001101_0010100100000000"; -- -0.3796820044517517
	pesos_i(8530) := b"1111111111111111_1111111111111111_1000010110001011_0110110010000000"; -- -0.47834131121635437
	pesos_i(8531) := b"0000000000000000_0000000000000000_0011010001101101_1011010000000000"; -- 0.20479893684387207
	pesos_i(8532) := b"0000000000000000_0000000000000000_0110011010101000_0000111110000000"; -- 0.401001900434494
	pesos_i(8533) := b"1111111111111111_1111111111111111_1011001001000010_1000101000000000"; -- -0.303672194480896
	pesos_i(8534) := b"1111111111111111_1111111111111111_1110111001001101_1011011101100000"; -- -0.06912664324045181
	pesos_i(8535) := b"0000000000000000_0000000000000000_0010101010101010_0010100101000000"; -- 0.16665895283222198
	pesos_i(8536) := b"1111111111111111_1111111111111111_1000100111001000_0000001000000000"; -- -0.46179187297821045
	pesos_i(8537) := b"0000000000000000_0000000000000000_0010011110110100_0000111011000000"; -- 0.15509121119976044
	pesos_i(8538) := b"0000000000000000_0000000000000000_0001011100011000_0100111110100000"; -- 0.09021470695734024
	pesos_i(8539) := b"1111111111111111_1111111111111111_1101010000111011_0011100110000000"; -- -0.17097130417823792
	pesos_i(8540) := b"0000000000000000_0000000000000000_0011101111101011_0010111000000000"; -- 0.23405730724334717
	pesos_i(8541) := b"1111111111111111_1111111111111111_1100010111100100_0100111000000000"; -- -0.22698509693145752
	pesos_i(8542) := b"0000000000000000_0000000000000000_0010010110111010_1010010011000000"; -- 0.14737920463085175
	pesos_i(8543) := b"1111111111111111_1111111111111111_0110100110001111_1001101100000000"; -- -0.5876525044441223
	pesos_i(8544) := b"1111111111111111_1111111111111111_1101010011111000_0001110001000000"; -- -0.1680891364812851
	pesos_i(8545) := b"1111111111111111_1111111111111111_1000110000111110_0011010010000000"; -- -0.4521758258342743
	pesos_i(8546) := b"1111111111111111_1111111111111111_1101001001111110_1100001010000000"; -- -0.1777532994747162
	pesos_i(8547) := b"0000000000000000_0000000000000000_0011011001010000_1011011111000000"; -- 0.21216915547847748
	pesos_i(8548) := b"0000000000000000_0000000000000000_0010110110010101_1111110010000000"; -- 0.1780698597431183
	pesos_i(8549) := b"0000000000000000_0000000000000000_0100100110100101_0000011110000000"; -- 0.2876743972301483
	pesos_i(8550) := b"1111111111111111_1111111111111111_1111110100100000_1111000000111000"; -- -0.011216150596737862
	pesos_i(8551) := b"1111111111111111_1111111111111111_1101000111010000_0001111001000000"; -- -0.18041811883449554
	pesos_i(8552) := b"0000000000000000_0000000000000000_0100111011111000_0101011000000000"; -- 0.3084768056869507
	pesos_i(8553) := b"0000000000000000_0000000000000000_0110100000100100_0011011110000000"; -- 0.40680262446403503
	pesos_i(8554) := b"1111111111111111_1111111111111111_0101110011111010_1111101100000000"; -- -0.6367953419685364
	pesos_i(8555) := b"0000000000000000_0000000000000000_0001110101111111_1111111101100000"; -- 0.11523433774709702
	pesos_i(8556) := b"1111111111111111_1111111111111111_0111010000101011_0111010000000000"; -- -0.5462119579315186
	pesos_i(8557) := b"0000000000000000_0000000000000000_0110110011111100_0010100100000000"; -- 0.4257226586341858
	pesos_i(8558) := b"0000000000000000_0000000000000000_0100100100111111_0100111000000000"; -- 0.28612220287323
	pesos_i(8559) := b"1111111111111111_1111111111111111_0111111001001001_0110010000000000"; -- -0.50669264793396
	pesos_i(8560) := b"1111111111111111_1111111111111111_1101010100101010_1000001010000000"; -- -0.1673201024532318
	pesos_i(8561) := b"1111111111111111_1111111111111111_1101100110101110_1001110001000000"; -- -0.14967940747737885
	pesos_i(8562) := b"1111111111111111_1111111111111111_1000101100111010_0010011110000000"; -- -0.45614388585090637
	pesos_i(8563) := b"0000000000000000_0000000000000000_0010011010000010_1000000100000000"; -- 0.15042883157730103
	pesos_i(8564) := b"0000000000000000_0000000000000000_0010001000111010_1011001101000000"; -- 0.133708193898201
	pesos_i(8565) := b"0000000000000000_0000000000000000_0011000000110100_1001011101000000"; -- 0.18830247223377228
	pesos_i(8566) := b"1111111111111111_1111111111111111_1111111111100110_1010000101000101"; -- -0.00038711607339791954
	pesos_i(8567) := b"0000000000000000_0000000000000000_0000001100000110_0110101101110100"; -- 0.01181670743972063
	pesos_i(8568) := b"0000000000000000_0000000000000000_0001101011001101_0010011010000000"; -- 0.10469284653663635
	pesos_i(8569) := b"1111111111111111_1111111111111111_1000110111011000_1101111110000000"; -- -0.4459095299243927
	pesos_i(8570) := b"0000000000000000_0000000000000000_0010101001101101_1011000110000000"; -- 0.16573628783226013
	pesos_i(8571) := b"1111111111111111_1111111111111111_1011101000110100_0011001100000000"; -- -0.27264100313186646
	pesos_i(8572) := b"1111111111111111_1111111111111111_0111110011111111_0000101100000000"; -- -0.51173335313797
	pesos_i(8573) := b"1111111111111111_1111111111111111_1110011100111100_1011101000000000"; -- -0.09672963619232178
	pesos_i(8574) := b"1111111111111111_1111111111111111_0110111001001101_0011011000000000"; -- -0.5691343545913696
	pesos_i(8575) := b"1111111111111111_1111111111111111_1110101101000100_0101101100000000"; -- -0.08098822832107544
	pesos_i(8576) := b"0000000000000000_0000000000000000_0110101101001110_0101010100000000"; -- 0.4191640019416809
	pesos_i(8577) := b"0000000000000000_0000000000000000_0000010100000111_0010101000100000"; -- 0.019640572369098663
	pesos_i(8578) := b"0000000000000000_0000000000000000_0000000101000111_0010011011110000"; -- 0.004991944879293442
	pesos_i(8579) := b"1111111111111111_1111111111111111_0101111000010101_0011001000000000"; -- -0.6324890851974487
	pesos_i(8580) := b"0000000000000000_0000000000000000_0110111010000010_1001000010000000"; -- 0.43167975544929504
	pesos_i(8581) := b"0000000000000000_0000000000000000_0010010011110110_1011111001000000"; -- 0.14439000189304352
	pesos_i(8582) := b"0000000000000000_0000000000000000_0111100011001110_0110110000000000"; -- 0.47189974784851074
	pesos_i(8583) := b"0000000000000000_0000000000000000_0010101101011100_1110101110000000"; -- 0.1693865954875946
	pesos_i(8584) := b"1111111111111111_1111111111111111_0110010100100111_1011100100000000"; -- -0.604862630367279
	pesos_i(8585) := b"1111111111111111_1111111111111111_1100001011101010_1110000001000000"; -- -0.23860357701778412
	pesos_i(8586) := b"0000000000000000_0000000000000000_0000100110111101_1101101101010000"; -- 0.0380532331764698
	pesos_i(8587) := b"0000000000000000_0000000000000000_0011010011010110_0011111111000000"; -- 0.20639418065547943
	pesos_i(8588) := b"1111111111111111_1111111111111111_1101111010111111_0101110011000000"; -- -0.12989254295825958
	pesos_i(8589) := b"0000000000000000_0000000000000000_0101110011110101_0000000110000000"; -- 0.36311349272727966
	pesos_i(8590) := b"1111111111111111_1111111111111111_1001100001111101_1011111100000000"; -- -0.4043312668800354
	pesos_i(8591) := b"0000000000000000_0000000000000000_0010111010100010_1000000100000000"; -- 0.18216711282730103
	pesos_i(8592) := b"1111111111111111_1111111111111111_1101101011010101_0011001010000000"; -- -0.14518436789512634
	pesos_i(8593) := b"1111111111111111_1111111111111111_1000100001111010_0011101100000000"; -- -0.46688491106033325
	pesos_i(8594) := b"1111111111111111_1111111111111111_1100001011110001_0100111000000000"; -- -0.23850548267364502
	pesos_i(8595) := b"0000000000000000_0000000000000000_0010010101000110_0111101000000000"; -- 0.1456066370010376
	pesos_i(8596) := b"1111111111111111_1111111111111111_0100001001001100_1001110100000000"; -- -0.7410184741020203
	pesos_i(8597) := b"0000000000000000_0000000000000000_0111111001000111_1100000010000000"; -- 0.49328234791755676
	pesos_i(8598) := b"0000000000000000_0000000000000000_0011011101000011_0110000010000000"; -- 0.21587184071540833
	pesos_i(8599) := b"1111111111111111_1111111111111110_1101010101101000_1010010000000000"; -- -1.1663720607757568
	pesos_i(8600) := b"1111111111111111_1111111111111111_1100001001110110_0110010100000000"; -- -0.24038094282150269
	pesos_i(8601) := b"1111111111111111_1111111111111111_1011010101011101_1100001000000000"; -- -0.2915381193161011
	pesos_i(8602) := b"0000000000000000_0000000000000000_0001111000100101_0110110001000000"; -- 0.11775852739810944
	pesos_i(8603) := b"0000000000000000_0000000000000000_0101000000000001_0101010100000000"; -- 0.3125203251838684
	pesos_i(8604) := b"0000000000000000_0000000000000000_0001000000110100_0111001000000000"; -- 0.0633002519607544
	pesos_i(8605) := b"0000000000000000_0000000000000000_0001000001000011_0100000100000000"; -- 0.0635262131690979
	pesos_i(8606) := b"1111111111111111_1111111111111111_0111111111011010_1010101100000000"; -- -0.5005696415901184
	pesos_i(8607) := b"1111111111111111_1111111111111111_1111011110100100_0011110011000000"; -- -0.032650187611579895
	pesos_i(8608) := b"0000000000000000_0000000000000000_0100001110101011_0010100000000000"; -- 0.2643303871154785
	pesos_i(8609) := b"1111111111111111_1111111111111111_1010111111111000_1101011000000000"; -- -0.31260931491851807
	pesos_i(8610) := b"0000000000000000_0000000000000000_0000011101000001_1001011110011000"; -- 0.02834460698068142
	pesos_i(8611) := b"0000000000000000_0000000000000000_0010011110010110_0100100000000000"; -- 0.15463685989379883
	pesos_i(8612) := b"0000000000000000_0000000000000000_0100000000100001_1011101110000000"; -- 0.2505147159099579
	pesos_i(8613) := b"0000000000000000_0000000000000000_0111010001110110_1000011110000000"; -- 0.45493361353874207
	pesos_i(8614) := b"1111111111111111_1111111111111111_1100101110100001_0111110100000000"; -- -0.20456713438034058
	pesos_i(8615) := b"0000000000000000_0000000000000000_0010001001010110_1011001100000000"; -- 0.1341354250907898
	pesos_i(8616) := b"1111111111111111_1111111111111111_1000110111100010_0100011000000000"; -- -0.4457660913467407
	pesos_i(8617) := b"1111111111111111_1111111111111111_1101111010010011_1111110101000000"; -- -0.13055436313152313
	pesos_i(8618) := b"0000000000000000_0000000000000000_0101010110101101_0010000010000000"; -- 0.3346729576587677
	pesos_i(8619) := b"1111111111111111_1111111111111111_1101101100111111_1010010110000000"; -- -0.14356008172035217
	pesos_i(8620) := b"0000000000000000_0000000000000000_0010011110010011_0000000110000000"; -- 0.15458688139915466
	pesos_i(8621) := b"1111111111111111_1111111111111111_1010101101000110_1010011010000000"; -- -0.3309532105922699
	pesos_i(8622) := b"1111111111111111_1111111111111111_1110100001011111_0100000010100000"; -- -0.09229656308889389
	pesos_i(8623) := b"0000000000000000_0000000000000000_1010011011010101_1100010000000000"; -- 0.6516993045806885
	pesos_i(8624) := b"1111111111111111_1111111111111111_1011000101010101_0011001100000000"; -- -0.30729371309280396
	pesos_i(8625) := b"1111111111111111_1111111111111111_1011111010101001_0101001010000000"; -- -0.25522884726524353
	pesos_i(8626) := b"1111111111111111_1111111111111111_1101110011101111_0111011100000000"; -- -0.13697105646133423
	pesos_i(8627) := b"1111111111111111_1111111111111111_0110101000010011_1001111100000000"; -- -0.5856381058692932
	pesos_i(8628) := b"0000000000000000_0000000000000000_0100100111101001_0000100000000000"; -- 0.2887120246887207
	pesos_i(8629) := b"0000000000000000_0000000000000000_0001110010001000_0101010000100000"; -- 0.11145520955324173
	pesos_i(8630) := b"1111111111111111_1111111111111111_1000100110001110_1110010000000000"; -- -0.4626634120941162
	pesos_i(8631) := b"0000000000000000_0000000000000000_0100110110100111_1110111100000000"; -- 0.3033437132835388
	pesos_i(8632) := b"1111111111111111_1111111111111111_1101010000100010_0001000010000000"; -- -0.1713552176952362
	pesos_i(8633) := b"0000000000000000_0000000000000000_0110100000000001_1101001000000000"; -- 0.40627777576446533
	pesos_i(8634) := b"0000000000000000_0000000000000000_0100010000000011_0001000110000000"; -- 0.26567181944847107
	pesos_i(8635) := b"0000000000000000_0000000000000000_0010100110110010_0111010110000000"; -- 0.1628793179988861
	pesos_i(8636) := b"1111111111111111_1111111111111111_1010001100001010_1110101000000000"; -- -0.36311471462249756
	pesos_i(8637) := b"1111111111111111_1111111111111111_1000111010011111_1100101010000000"; -- -0.4428742825984955
	pesos_i(8638) := b"1111111111111111_1111111111111110_1111100001110101_1100001000000000"; -- -1.029453158378601
	pesos_i(8639) := b"0000000000000000_0000000000000000_0011100101111000_0001001001000000"; -- 0.22448839247226715
	pesos_i(8640) := b"1111111111111111_1111111111111111_1110110000010001_1001001010000000"; -- -0.0778568685054779
	pesos_i(8641) := b"0000000000000000_0000000000000000_0011000101001000_0101100000000000"; -- 0.19251012802124023
	pesos_i(8642) := b"0000000000000000_0000000000000000_0101110011000000_0111100000000000"; -- 0.36231184005737305
	pesos_i(8643) := b"1111111111111111_1111111111111111_1100000000010101_0000010010000000"; -- -0.249679297208786
	pesos_i(8644) := b"0000000000000000_0000000000000000_0101011000101010_1001110010000000"; -- 0.33658769726753235
	pesos_i(8645) := b"0000000000000000_0000000000000000_0000011111011110_0111010110011000"; -- 0.030738210305571556
	pesos_i(8646) := b"1111111111111111_1111111111111111_0101000001100110_1111010100000000"; -- -0.685929000377655
	pesos_i(8647) := b"1111111111111111_1111111111111111_1110010001000001_0100001010000000"; -- -0.10837921500205994
	pesos_i(8648) := b"0000000000000000_0000000000000000_0010010001010001_0010100101000000"; -- 0.14186342060565948
	pesos_i(8649) := b"1111111111111111_1111111111111111_1110001011110011_0000001101000000"; -- -0.11347942054271698
	pesos_i(8650) := b"0000000000000000_0000000000000000_0100001111110110_1011001000000000"; -- 0.265483021736145
	pesos_i(8651) := b"1111111111111111_1111111111111111_1101110111111110_1101101101000000"; -- -0.132829949259758
	pesos_i(8652) := b"1111111111111111_1111111111111111_0000011101111100_1111110000000000"; -- -0.9707491397857666
	pesos_i(8653) := b"1111111111111111_1111111111111111_1110100100010010_0100001010000000"; -- -0.08956512808799744
	pesos_i(8654) := b"0000000000000000_0000000000000000_0001111101000010_0111101111100000"; -- 0.12210821360349655
	pesos_i(8655) := b"0000000000000000_0000000000000000_0000111010010011_1000011000000000"; -- 0.0569385290145874
	pesos_i(8656) := b"0000000000000000_0000000000000000_0001110111010011_1100010100100000"; -- 0.11651260405778885
	pesos_i(8657) := b"1111111111111111_1111111111111111_1101110001101011_0100011011000000"; -- -0.13898809254169464
	pesos_i(8658) := b"1111111111111111_1111111111111111_1010111001110011_1100110110000000"; -- -0.31854549050331116
	pesos_i(8659) := b"0000000000000000_0000000000000000_0101110011101001_1111101100000000"; -- 0.3629452586174011
	pesos_i(8660) := b"1111111111111111_1111111111111111_1000001011010000_1110011000000000"; -- -0.48899996280670166
	pesos_i(8661) := b"0000000000000000_0000000000000000_0101101001010111_1011011000000000"; -- 0.3529008626937866
	pesos_i(8662) := b"0000000000000000_0000000000000000_0011111000111100_0001100111000000"; -- 0.24310456216335297
	pesos_i(8663) := b"1111111111111111_1111111111111111_0110010111110000_0011110000000000"; -- -0.6018030643463135
	pesos_i(8664) := b"0000000000000000_0000000000000000_0000101000010100_0111011001100000"; -- 0.03937473148107529
	pesos_i(8665) := b"1111111111111111_1111111111111111_1101101010101111_1001111100000000"; -- -0.1457577347755432
	pesos_i(8666) := b"1111111111111111_1111111111111111_0101011011000000_0011111100000000"; -- -0.6611290574073792
	pesos_i(8667) := b"0000000000000000_0000000000000000_0110010110011110_0000011000000000"; -- 0.39694249629974365
	pesos_i(8668) := b"1111111111111111_1111111111111111_1101111001110110_0110101110000000"; -- -0.13100555539131165
	pesos_i(8669) := b"0000000000000000_0000000000000000_0010011010001110_0100111111000000"; -- 0.15060900151729584
	pesos_i(8670) := b"0000000000000000_0000000000000000_0100001110100111_1101110010000000"; -- 0.2642801105976105
	pesos_i(8671) := b"1111111111111111_1111111111111111_0111110001011101_0111110000000000"; -- -0.5141985416412354
	pesos_i(8672) := b"0000000000000000_0000000000000000_0000101000101000_1100101011010000"; -- 0.03968494012951851
	pesos_i(8673) := b"0000000000000000_0000000000000000_0101011111001000_1110010100000000"; -- 0.34290915727615356
	pesos_i(8674) := b"1111111111111111_1111111111111111_1111000111001000_1101000111110000"; -- -0.055529478937387466
	pesos_i(8675) := b"0000000000000000_0000000000000000_0011001111101110_0010000110000000"; -- 0.20285233855247498
	pesos_i(8676) := b"1111111111111111_1111111111111111_0111010100101000_0111001100000000"; -- -0.5423515439033508
	pesos_i(8677) := b"1111111111111111_1111111111111111_1110000000110000_1000000011000000"; -- -0.12425990402698517
	pesos_i(8678) := b"1111111111111111_1111111111111111_1100100111100010_0001000000000000"; -- -0.2113943099975586
	pesos_i(8679) := b"1111111111111111_1111111111111111_0101111011100111_0010100000000000"; -- -0.6292853355407715
	pesos_i(8680) := b"0000000000000000_0000000000000000_0100110101001100_0001010000000000"; -- 0.3019421100616455
	pesos_i(8681) := b"1111111111111111_1111111111111111_1011110001111011_1011001000000000"; -- -0.2637375593185425
	pesos_i(8682) := b"1111111111111111_1111111111111111_1111111001100000_1100010000011010"; -- -0.0063359676860272884
	pesos_i(8683) := b"0000000000000000_0000000000000000_0111000001100010_0100000010000000"; -- 0.438999205827713
	pesos_i(8684) := b"0000000000000000_0000000000000000_0100110000000101_1010101100000000"; -- 0.2969614863395691
	pesos_i(8685) := b"1111111111111111_1111111111111111_0101101101001100_1100100100000000"; -- -0.6433596014976501
	pesos_i(8686) := b"0000000000000000_0000000000000000_0011001111010111_1011111100000000"; -- 0.2025107741355896
	pesos_i(8687) := b"1111111111111111_1111111111111111_0101100010001101_0110000000000000"; -- -0.6540927886962891
	pesos_i(8688) := b"0000000000000000_0000000000000000_0011010101010011_1001011010000000"; -- 0.2083066999912262
	pesos_i(8689) := b"0000000000000000_0000000000000000_1001111000110010_1111000100000000"; -- 0.6179648041725159
	pesos_i(8690) := b"1111111111111111_1111111111111111_0110000010001110_0101110000000000"; -- -0.6228277683258057
	pesos_i(8691) := b"1111111111111111_1111111111111111_0011001100000110_1101101100000000"; -- -0.8006766438484192
	pesos_i(8692) := b"1111111111111111_1111111111111111_1100011110111001_0001110000000000"; -- -0.2198317050933838
	pesos_i(8693) := b"0000000000000000_0000000000000000_0011111010111111_1110001101000000"; -- 0.2451154738664627
	pesos_i(8694) := b"1111111111111111_1111111111111111_0111011100111101_1100000000000000"; -- -0.5342140197753906
	pesos_i(8695) := b"0000000000000000_0000000000000000_0001001000100110_1110101010000000"; -- 0.07090631127357483
	pesos_i(8696) := b"0000000000000000_0000000000000000_0101011110100000_0101101000000000"; -- 0.3422905206680298
	pesos_i(8697) := b"1111111111111111_1111111111111111_1110010101001010_1101010110000000"; -- -0.10432687401771545
	pesos_i(8698) := b"0000000000000000_0000000000000000_0000101100110110_1111010001110000"; -- 0.043807294219732285
	pesos_i(8699) := b"1111111111111111_1111111111111111_1100111111011010_0010100011000000"; -- -0.1880774050951004
	pesos_i(8700) := b"0000000000000000_0000000000000000_0010110101000010_0111001011000000"; -- 0.17679516971111298
	pesos_i(8701) := b"0000000000000000_0000000000000000_0101001111111000_0101010100000000"; -- 0.3280079960823059
	pesos_i(8702) := b"1111111111111111_1111111111111111_0100110010001011_1001001100000000"; -- -0.7009952664375305
	pesos_i(8703) := b"0000000000000000_0000000000000000_0101111001010001_1000100010000000"; -- 0.36843159794807434
	pesos_i(8704) := b"1111111111111111_1111111111111111_1110001010010101_0001111010100000"; -- -0.11491211503744125
	pesos_i(8705) := b"1111111111111111_1111111111111111_0110101001010001_1000110000000000"; -- -0.584693193435669
	pesos_i(8706) := b"1111111111111111_1111111111111111_0000000100101110_1001000100000000"; -- -0.9953832030296326
	pesos_i(8707) := b"0000000000000000_0000000000000000_1101011101111111_1000110100000000"; -- 0.8417900204658508
	pesos_i(8708) := b"0000000000000000_0000000000000000_1001110101111100_1011011000000000"; -- 0.6151841878890991
	pesos_i(8709) := b"0000000000000000_0000000000000000_0001110101100010_0101100100100000"; -- 0.1147819235920906
	pesos_i(8710) := b"1111111111111111_1111111111111111_1101001100110111_1100111011000000"; -- -0.1749296933412552
	pesos_i(8711) := b"0000000000000000_0000000000000000_0011100001101100_0011100101000000"; -- 0.2204013615846634
	pesos_i(8712) := b"0000000000000000_0000000000000000_0110100111111100_1000000000000000"; -- 0.41400909423828125
	pesos_i(8713) := b"1111111111111111_1111111111111111_0110101011110000_1110010100000000"; -- -0.5822617411613464
	pesos_i(8714) := b"1111111111111111_1111111111111111_1100101100001100_1111001111000000"; -- -0.206833615899086
	pesos_i(8715) := b"1111111111111111_1111111111111111_1110111000111001_0101000010100000"; -- -0.06943794339895248
	pesos_i(8716) := b"0000000000000000_0000000000000000_0000001010101100_0000000110100000"; -- 0.01043710857629776
	pesos_i(8717) := b"0000000000000000_0000000000000000_0010100111111100_1111000101000000"; -- 0.16401584446430206
	pesos_i(8718) := b"1111111111111111_1111111111111111_1101010110000100_0111001000000000"; -- -0.1659477949142456
	pesos_i(8719) := b"0000000000000000_0000000000000000_0010000101101001_0111111011000000"; -- 0.13051597774028778
	pesos_i(8720) := b"0000000000000000_0000000000000000_0001101001110110_0101011001100000"; -- 0.10336818546056747
	pesos_i(8721) := b"0000000000000000_0000000000000000_0100000110010010_1010001010000000"; -- 0.256143718957901
	pesos_i(8722) := b"1111111111111111_1111111111111111_1110111011000100_1111110111000000"; -- -0.06730665266513824
	pesos_i(8723) := b"0000000000000000_0000000000000000_0101000011011101_1011000010000000"; -- 0.31588271260261536
	pesos_i(8724) := b"1111111111111111_1111111111111111_1001001111100010_0001101110000000"; -- -0.4223311245441437
	pesos_i(8725) := b"1111111111111111_1111111111111111_1110111111111010_0001101001000000"; -- -0.06258998811244965
	pesos_i(8726) := b"0000000000000000_0000000000000000_0110100011111010_1100110010000000"; -- 0.41007688641548157
	pesos_i(8727) := b"1111111111111111_1111111111111111_1111001001101000_0100000000110000"; -- -0.05309676006436348
	pesos_i(8728) := b"1111111111111111_1111111111111111_0111100111101011_0110111000000000"; -- -0.5237513780593872
	pesos_i(8729) := b"1111111111111111_1111111111111111_1111111100010011_1101100101110001"; -- -0.0036033724900335073
	pesos_i(8730) := b"0000000000000000_0000000000000000_0011000011000011_1111000100000000"; -- 0.19048982858657837
	pesos_i(8731) := b"0000000000000000_0000000000000000_0000111011011101_0011101100110000"; -- 0.05806322023272514
	pesos_i(8732) := b"1111111111111111_1111111111111111_1101111111010110_0010100001000000"; -- -0.1256384700536728
	pesos_i(8733) := b"1111111111111111_1111111111111111_1111101001101011_1010101001001000"; -- -0.02179466001689434
	pesos_i(8734) := b"0000000000000000_0000000000000000_0101010000011101_1000001010000000"; -- 0.3285752832889557
	pesos_i(8735) := b"0000000000000000_0000000000000000_0000110010100100_1011010001010000"; -- 0.04938818886876106
	pesos_i(8736) := b"1111111111111111_1111111111111111_1100110110101101_0110011010000000"; -- -0.19657287001609802
	pesos_i(8737) := b"0000000000000000_0000000000000000_0010110010111100_0101011001000000"; -- 0.17474879324436188
	pesos_i(8738) := b"0000000000000000_0000000000000000_0000101101111010_0000111000100000"; -- 0.04483116418123245
	pesos_i(8739) := b"1111111111111111_1111111111111111_0110101001000111_1011000000000000"; -- -0.584843635559082
	pesos_i(8740) := b"0000000000000000_0000000000000000_0101100100011001_1011001110000000"; -- 0.3480484187602997
	pesos_i(8741) := b"1111111111111111_1111111111111111_0111000011110000_1000000100000000"; -- -0.558830201625824
	pesos_i(8742) := b"1111111111111111_1111111111111111_1100111111111110_0001011111000000"; -- -0.18752910196781158
	pesos_i(8743) := b"1111111111111111_1111111111111111_0111011000000000_0110001100000000"; -- -0.5390565991401672
	pesos_i(8744) := b"0000000000000000_0000000000000000_0001100001000100_0001001010100000"; -- 0.09478870779275894
	pesos_i(8745) := b"0000000000000000_0000000000000000_0101011011111110_1100011100000000"; -- 0.3398250937461853
	pesos_i(8746) := b"1111111111111111_1111111111111111_1101010111110011_1010011000000000"; -- -0.16425096988677979
	pesos_i(8747) := b"0000000000000000_0000000000000000_0000100100011001_0100100011010000"; -- 0.03554205968976021
	pesos_i(8748) := b"1111111111111111_1111111111111111_0000000011110101_0101110000000000"; -- -0.9962561130523682
	pesos_i(8749) := b"0000000000000000_0000000000000000_0101011001001110_0111010110000000"; -- 0.3371346890926361
	pesos_i(8750) := b"0000000000000000_0000000000000000_0010001001101000_0100100100000000"; -- 0.1344037652015686
	pesos_i(8751) := b"0000000000000000_0000000000000000_0010001001000001_0111100010000000"; -- 0.13381150364875793
	pesos_i(8752) := b"1111111111111111_1111111111111111_0001110000100111_0111101100000000"; -- -0.8900225758552551
	pesos_i(8753) := b"0000000000000000_0000000000000000_0100111000110101_0000110100000000"; -- 0.3054969906806946
	pesos_i(8754) := b"1111111111111111_1111111111111111_1100110000101001_0100111111000000"; -- -0.20249463617801666
	pesos_i(8755) := b"1111111111111111_1111111111111111_1001100010000111_1111000100000000"; -- -0.40417569875717163
	pesos_i(8756) := b"0000000000000000_0000000000000000_0101100010111001_1010000010000000"; -- 0.34658244252204895
	pesos_i(8757) := b"0000000000000000_0000000000000000_0010110011101110_0010000100000000"; -- 0.1755085587501526
	pesos_i(8758) := b"1111111111111111_1111111111111111_1110111010100110_1101001111100000"; -- -0.06776691228151321
	pesos_i(8759) := b"1111111111111111_1111111111111111_1110100110111101_0001100010100000"; -- -0.0869583711028099
	pesos_i(8760) := b"0000000000000000_0000000000000000_0011011111111110_0101011110000000"; -- 0.21872469782829285
	pesos_i(8761) := b"0000000000000000_0000000000000000_0001010100101100_1110100110100000"; -- 0.08271656185388565
	pesos_i(8762) := b"1111111111111111_1111111111111111_1000000011100010_0011011010000000"; -- -0.49654826521873474
	pesos_i(8763) := b"0000000000000000_0000000000000000_0011000111000100_1001111001000000"; -- 0.1944064050912857
	pesos_i(8764) := b"0000000000000000_0000000000000000_0100100000011100_0000110010000000"; -- 0.2816779911518097
	pesos_i(8765) := b"0000000000000000_0000000000000000_0110000110111001_1100101000000000"; -- 0.38174116611480713
	pesos_i(8766) := b"1111111111111111_1111111111111111_0101000100110010_0100000100000000"; -- -0.6828269362449646
	pesos_i(8767) := b"0000000000000000_0000000000000000_0001001001000011_0110010010100000"; -- 0.07134083658456802
	pesos_i(8768) := b"1111111111111111_1111111111111111_0001111000110000_0000111000000000"; -- -0.8820792436599731
	pesos_i(8769) := b"0000000000000000_0000000000000000_0100001001000111_1010011100000000"; -- 0.258905827999115
	pesos_i(8770) := b"0000000000000000_0000000000000000_0000011110111100_1100111100111000"; -- 0.03022475354373455
	pesos_i(8771) := b"0000000000000000_0000000000000000_0001111011101110_1001001000000000"; -- 0.12082779407501221
	pesos_i(8772) := b"1111111111111111_1111111111111111_1010101101001101_0010001110000000"; -- -0.330854207277298
	pesos_i(8773) := b"1111111111111111_1111111111111111_1101111111100011_1000000010000000"; -- -0.12543484568595886
	pesos_i(8774) := b"1111111111111111_1111111111111111_0111111011011111_1001101100000000"; -- -0.5044005513191223
	pesos_i(8775) := b"1111111111111111_1111111111111111_1010011011111110_1101011010000000"; -- -0.3476739823818207
	pesos_i(8776) := b"0000000000000000_0000000000000000_0010010111111001_0100001001000000"; -- 0.14833463728427887
	pesos_i(8777) := b"1111111111111111_1111111111111111_1010001000010101_1010011100000000"; -- -0.36685711145401
	pesos_i(8778) := b"1111111111111111_1111111111111111_1111000101010001_0000110100100000"; -- -0.05735700577497482
	pesos_i(8779) := b"0000000000000000_0000000000000000_0100011010001111_1001001000000000"; -- 0.2756282091140747
	pesos_i(8780) := b"0000000000000000_0000000000000000_0001111000010011_0101011011100000"; -- 0.11748259514570236
	pesos_i(8781) := b"0000000000000000_0000000000000000_0100111111000000_1100001110000000"; -- 0.3115350902080536
	pesos_i(8782) := b"0000000000000000_0000000000000000_0000110000011000_0001101111000000"; -- 0.04724286496639252
	pesos_i(8783) := b"0000000000000000_0000000000000000_0010110111000110_0100110000000000"; -- 0.17880702018737793
	pesos_i(8784) := b"1111111111111111_1111111111111111_1111100000111000_1110010000101000"; -- -0.030381908640265465
	pesos_i(8785) := b"0000000000000000_0000000000000000_0101110101011111_1001101100000000"; -- 0.3647400736808777
	pesos_i(8786) := b"1111111111111111_1111111111111111_1000011011100001_0011001110000000"; -- -0.47312620282173157
	pesos_i(8787) := b"0000000000000000_0000000000000000_0000101100010000_1011100100100000"; -- 0.043223924934864044
	pesos_i(8788) := b"0000000000000000_0000000000000000_0001101011111110_0100101001000000"; -- 0.10544265806674957
	pesos_i(8789) := b"1111111111111111_1111111111111111_1101111011111011_0000101100000000"; -- -0.12898188829421997
	pesos_i(8790) := b"1111111111111111_1111111111111111_1111110011000111_0010011110001000"; -- -0.012586144730448723
	pesos_i(8791) := b"1111111111111111_1111111111111111_1011111110101011_0000000000000000"; -- -0.2512969970703125
	pesos_i(8792) := b"1111111111111111_1111111111111111_1011101101000011_0010111000000000"; -- -0.26850616931915283
	pesos_i(8793) := b"0000000000000000_0000000000000000_0000111000101100_1100100000100000"; -- 0.055370815098285675
	pesos_i(8794) := b"0000000000000000_0000000000000000_0001100001000000_1100001011100000"; -- 0.0947381779551506
	pesos_i(8795) := b"0000000000000000_0000000000000000_0010101010101010_0010010011000000"; -- 0.1666586846113205
	pesos_i(8796) := b"1111111111111111_1111111111111111_1110000100100101_0100100010000000"; -- -0.12052485346794128
	pesos_i(8797) := b"1111111111111111_1111111111111111_1011110001000101_1100111010000000"; -- -0.2645598351955414
	pesos_i(8798) := b"1111111111111111_1111111111111111_1001110101001101_1011111000000000"; -- -0.3855324983596802
	pesos_i(8799) := b"0000000000000000_0000000000000000_0000000001011100_1010101101101100"; -- 0.0014140261337161064
	pesos_i(8800) := b"0000000000000000_0000000000000000_0100101110000001_0110111000000000"; -- 0.2949436902999878
	pesos_i(8801) := b"1111111111111111_1111111111111111_1111111010000111_1001001011000010"; -- -0.005743816029280424
	pesos_i(8802) := b"1111111111111111_1111111111111111_1111010100001001_1001000001010000"; -- -0.04282281920313835
	pesos_i(8803) := b"1111111111111111_1111111111111111_1111100111111010_0100111111000000"; -- -0.023524299263954163
	pesos_i(8804) := b"0000000000000000_0000000000000000_0000000001110000_0010111011101110"; -- 0.0017117816023528576
	pesos_i(8805) := b"1111111111111111_1111111111111111_0011000010001001_0011001000000000"; -- -0.8104065656661987
	pesos_i(8806) := b"0000000000000000_0000000000000000_0001111100001001_0110000001100000"; -- 0.12123682349920273
	pesos_i(8807) := b"1111111111111111_1111111111111111_1111010110011100_0000110010010000"; -- -0.04058763012290001
	pesos_i(8808) := b"0000000000000000_0000000000000000_0010100110010110_0101110010000000"; -- 0.16245058178901672
	pesos_i(8809) := b"1111111111111111_1111111111111111_0011010000100100_0010110000000000"; -- -0.7963230609893799
	pesos_i(8810) := b"0000000000000000_0000000000000000_0011001000101001_0101011011000000"; -- 0.19594328105449677
	pesos_i(8811) := b"0000000000000000_0000000000000000_0011100111000011_1011001100000000"; -- 0.2256423830986023
	pesos_i(8812) := b"1111111111111111_1111111111111111_0111111011010000_1011111100000000"; -- -0.5046272873878479
	pesos_i(8813) := b"1111111111111111_1111111111111111_1011110111000001_0000001110000000"; -- -0.2587735950946808
	pesos_i(8814) := b"1111111111111111_1111111111111111_1111101101110100_0101110000000000"; -- -0.017755746841430664
	pesos_i(8815) := b"0000000000000000_0000000000000000_0001100100010111_0001111011000000"; -- 0.09800903499126434
	pesos_i(8816) := b"0000000000000000_0000000000000000_0000111011011111_1101001101000000"; -- 0.0581028014421463
	pesos_i(8817) := b"1111111111111111_1111111111111111_1101100011011011_1000010100000000"; -- -0.15290039777755737
	pesos_i(8818) := b"1111111111111111_1111111111111111_1111101111000000_0110110101011000"; -- -0.01659504510462284
	pesos_i(8819) := b"0000000000000000_0000000000000000_0100111001100010_0001010000000000"; -- 0.3061840534210205
	pesos_i(8820) := b"1111111111111111_1111111111111111_1101100000000100_0111001000000000"; -- -0.1561821699142456
	pesos_i(8821) := b"1111111111111111_1111111111111111_1000101110100110_0110100110000000"; -- -0.4544920027256012
	pesos_i(8822) := b"1111111111111111_1111111111111111_1110010001010011_1101010111000000"; -- -0.10809578001499176
	pesos_i(8823) := b"1111111111111111_1111111111111111_1101100010010010_0111011100000000"; -- -0.15401512384414673
	pesos_i(8824) := b"0000000000000000_0000000000000000_0010001101111001_1000010000000000"; -- 0.13857293128967285
	pesos_i(8825) := b"1111111111111111_1111111111111111_0010010001000111_0001111000000000"; -- -0.8582898378372192
	pesos_i(8826) := b"1111111111111111_1111111111111111_0111101000001000_0010110100000000"; -- -0.5233127474784851
	pesos_i(8827) := b"0000000000000000_0000000000000000_1000111101010101_1110001000000000"; -- 0.5599042177200317
	pesos_i(8828) := b"0000000000000000_0000000000000000_1001010110110100_0101101000000000"; -- 0.5847831964492798
	pesos_i(8829) := b"1111111111111111_1111111111111111_0111101100011000_0010010000000000"; -- -0.5191628932952881
	pesos_i(8830) := b"1111111111111111_1111111111111111_1000110011001011_1110011110000000"; -- -0.450013667345047
	pesos_i(8831) := b"1111111111111111_1111111111111111_0110111101110011_1100110000000000"; -- -0.5646393299102783
	pesos_i(8832) := b"1111111111111111_1111111111111111_0100011000110011_1100101000000000"; -- -0.7257722616195679
	pesos_i(8833) := b"1111111111111111_1111111111111111_0111000110111001_1110001100000000"; -- -0.5557573437690735
	pesos_i(8834) := b"0000000000000000_0000000000000000_0101011011101101_1101001000000000"; -- 0.33956634998321533
	pesos_i(8835) := b"1111111111111111_1111111111111111_1000111100101001_1101101000000000"; -- -0.44076764583587646
	pesos_i(8836) := b"0000000000000000_0000000000000000_0100100001000001_0100010000000000"; -- 0.2822458744049072
	pesos_i(8837) := b"0000000000000000_0000000000000000_1101110111010000_0001011100000000"; -- 0.8664564490318298
	pesos_i(8838) := b"0000000000000000_0000000000000000_0011100111110001_0000100010000000"; -- 0.2263341248035431
	pesos_i(8839) := b"1111111111111111_1111111111111111_1011100100111100_1101011000000000"; -- -0.27641546726226807
	pesos_i(8840) := b"1111111111111111_1111111111111111_1010000111110101_1100010010000000"; -- -0.36734363436698914
	pesos_i(8841) := b"1111111111111111_1111111111111111_1000100010111001_1000101100000000"; -- -0.4659188389778137
	pesos_i(8842) := b"0000000000000000_0000000000000000_0000000100101010_0110011011101000"; -- 0.0045532528311014175
	pesos_i(8843) := b"0000000000000000_0000000000000000_0101100101110011_0011111100000000"; -- 0.34941476583480835
	pesos_i(8844) := b"1111111111111111_1111111111111110_1111101000100111_0100100000000000"; -- -1.0228381156921387
	pesos_i(8845) := b"1111111111111111_1111111111111111_1101000100001000_1111000011000000"; -- -0.18345732986927032
	pesos_i(8846) := b"1111111111111111_1111111111111111_1100000101100110_1010010000000000"; -- -0.24452757835388184
	pesos_i(8847) := b"0000000000000000_0000000000000000_1010101010100001_0001101000000000"; -- 0.6665207147598267
	pesos_i(8848) := b"0000000000000000_0000000000000000_0001001110000101_1001100110100000"; -- 0.07625732570886612
	pesos_i(8849) := b"0000000000000000_0000000000000000_0011011001100000_1001101011000000"; -- 0.212411567568779
	pesos_i(8850) := b"1111111111111111_1111111111111111_0100001100110101_0111111100000000"; -- -0.737464964389801
	pesos_i(8851) := b"1111111111111111_1111111111111111_1100100111000101_0101111011000000"; -- -0.21183212101459503
	pesos_i(8852) := b"1111111111111111_1111111111111111_0110010111001100_0111101000000000"; -- -0.6023486852645874
	pesos_i(8853) := b"0000000000000000_0000000000000000_0101101101010111_0000101010000000"; -- 0.35679689049720764
	pesos_i(8854) := b"0000000000000000_0000000000000000_0100011010110111_0111001010000000"; -- 0.2762366831302643
	pesos_i(8855) := b"1111111111111111_1111111111111111_1111100001001000_0111101011100000"; -- -0.030144043266773224
	pesos_i(8856) := b"1111111111111111_1111111111111111_1011011101000000_0010010110000000"; -- -0.2841774523258209
	pesos_i(8857) := b"0000000000000000_0000000000000000_0010100110101101_1000000111000000"; -- 0.1628037542104721
	pesos_i(8858) := b"1111111111111111_1111111111111111_1111100001110000_1111010110100000"; -- -0.029526375234127045
	pesos_i(8859) := b"1111111111111111_1111111111111111_1010011000101010_0100111000000000"; -- -0.3509169816970825
	pesos_i(8860) := b"0000000000000000_0000000000000000_0100010010001010_1001011000000000"; -- 0.2677396535873413
	pesos_i(8861) := b"0000000000000000_0000000000000000_0001110101011101_0100101011100000"; -- 0.11470478028059006
	pesos_i(8862) := b"0000000000000000_0000000000000000_0100100101101101_1111111000000000"; -- 0.28683459758758545
	pesos_i(8863) := b"1111111111111111_1111111111111111_1000110110100110_1010101010000000"; -- -0.4466756284236908
	pesos_i(8864) := b"0000000000000000_0000000000000000_0011011111101101_1010011101000000"; -- 0.21847005188465118
	pesos_i(8865) := b"1111111111111111_1111111111111111_1111001100010011_0010001001110000"; -- -0.05048928037285805
	pesos_i(8866) := b"1111111111111111_1111111111111111_1001001110110010_0001011110000000"; -- -0.4230637848377228
	pesos_i(8867) := b"0000000000000000_0000000000000000_0010101000110110_0100110010000000"; -- 0.16489103436470032
	pesos_i(8868) := b"1111111111111111_1111111111111111_1100111111100100_1000101010000000"; -- -0.1879189908504486
	pesos_i(8869) := b"1111111111111111_1111111111111111_0111101101100101_0010100100000000"; -- -0.5179876685142517
	pesos_i(8870) := b"1111111111111111_1111111111111111_1111111101111100_1100111110010001"; -- -0.0020017882343381643
	pesos_i(8871) := b"1111111111111111_1111111111111111_1101011111100110_0010101011000000"; -- -0.15664418041706085
	pesos_i(8872) := b"1111111111111111_1111111111111111_1000001100100100_0101100000000000"; -- -0.48772668838500977
	pesos_i(8873) := b"0000000000000000_0000000000000000_0011111100011000_0110100010000000"; -- 0.24646618962287903
	pesos_i(8874) := b"1111111111111111_1111111111111111_0111110111001011_1010000100000000"; -- -0.5086116194725037
	pesos_i(8875) := b"0000000000000000_0000000000000000_0101110010100101_1000100110000000"; -- 0.3619008958339691
	pesos_i(8876) := b"0000000000000000_0000000000000000_0101100110001100_0100000100000000"; -- 0.3497963547706604
	pesos_i(8877) := b"1111111111111111_1111111111111111_1110010001001100_0100110111000000"; -- -0.10821069777011871
	pesos_i(8878) := b"1111111111111111_1111111111111111_0111111000011011_0000111100000000"; -- -0.5073996186256409
	pesos_i(8879) := b"0000000000000000_0000000000000000_0101011001110001_0100011100000000"; -- 0.33766597509384155
	pesos_i(8880) := b"1111111111111111_1111111111111111_1010101110011110_1101110010000000"; -- -0.329607218503952
	pesos_i(8881) := b"1111111111111111_1111111111111111_1101110010101011_1001010100000000"; -- -0.13800686597824097
	pesos_i(8882) := b"1111111111111111_1111111111111111_1010000011010001_0010001110000000"; -- -0.371808797121048
	pesos_i(8883) := b"0000000000000000_0000000000000000_0101011000110011_0111111100000000"; -- 0.336723268032074
	pesos_i(8884) := b"0000000000000000_0000000000000000_0101101000111000_1110001000000000"; -- 0.35243046283721924
	pesos_i(8885) := b"0000000000000000_0000000000000000_0010100101100100_1101111111000000"; -- 0.1616954654455185
	pesos_i(8886) := b"1111111111111111_1111111111111111_1100001101110111_0011001001000000"; -- -0.23646245896816254
	pesos_i(8887) := b"1111111111111111_1111111111111111_1001110111101011_0011011010000000"; -- -0.38312968611717224
	pesos_i(8888) := b"0000000000000000_0000000000000000_0011000001011010_0110110100000000"; -- 0.18887978792190552
	pesos_i(8889) := b"0000000000000000_0000000000000000_0101000111010100_0100111000000000"; -- 0.3196457624435425
	pesos_i(8890) := b"1111111111111111_1111111111111111_1110111010110010_0010000010100000"; -- -0.0675944909453392
	pesos_i(8891) := b"1111111111111111_1111111111111111_0101011010000000_1101001100000000"; -- -0.6620967984199524
	pesos_i(8892) := b"0000000000000000_0000000000000000_0011011100011011_0110011001000000"; -- 0.21526183187961578
	pesos_i(8893) := b"0000000000000000_0000000000000000_0001101000111011_1100100001000000"; -- 0.10247470438480377
	pesos_i(8894) := b"1111111111111111_1111111111111110_1010110010000101_1000010000000000"; -- -1.3260877132415771
	pesos_i(8895) := b"1111111111111111_1111111111111111_0011110100101011_1010000000000000"; -- -0.7610530853271484
	pesos_i(8896) := b"1111111111111111_1111111111111111_1001010110010011_1011000000000000"; -- -0.41571521759033203
	pesos_i(8897) := b"0000000000000000_0000000000000000_1000101011110101_1000110000000000"; -- 0.542809247970581
	pesos_i(8898) := b"0000000000000000_0000000000000000_0010110011110101_0111110101000000"; -- 0.17562086880207062
	pesos_i(8899) := b"0000000000000000_0000000000000000_0011110001001011_1000100000000000"; -- 0.23552751541137695
	pesos_i(8900) := b"0000000000000000_0000000000000000_0100101101111000_1100101000000000"; -- 0.29481184482574463
	pesos_i(8901) := b"0000000000000000_0000000000000000_0101110111101110_0111000110000000"; -- 0.366919606924057
	pesos_i(8902) := b"1111111111111111_1111111111111111_1000101111010001_0111101100000000"; -- -0.4538348317146301
	pesos_i(8903) := b"1111111111111111_1111111111111111_0111101010010101_0110100100000000"; -- -0.5211576819419861
	pesos_i(8904) := b"0000000000000000_0000000000000000_0001010100011101_0110101111000000"; -- 0.08248017728328705
	pesos_i(8905) := b"1111111111111111_1111111111111111_1111010110010010_0000100110110000"; -- -0.04074038937687874
	pesos_i(8906) := b"0000000000000000_0000000000000000_0100001110111001_0110101000000000"; -- 0.2645479440689087
	pesos_i(8907) := b"1111111111111111_1111111111111111_1000011000101111_1010001110000000"; -- -0.4758355915546417
	pesos_i(8908) := b"1111111111111111_1111111111111111_1001101000110100_0000000010000000"; -- -0.3976440131664276
	pesos_i(8909) := b"1111111111111111_1111111111111111_1110011011011011_1010100101000000"; -- -0.09821073710918427
	pesos_i(8910) := b"0000000000000000_0000000000000000_0001011101011000_1111000011000000"; -- 0.09120087325572968
	pesos_i(8911) := b"0000000000000000_0000000000000000_0001000101010111_0011001011000000"; -- 0.06773678958415985
	pesos_i(8912) := b"0000000000000000_0000000000000000_0111010000010011_1010111100000000"; -- 0.4534253478050232
	pesos_i(8913) := b"1111111111111111_1111111111111111_1010011011101111_1001010110000000"; -- -0.3479067385196686
	pesos_i(8914) := b"0000000000000000_0000000000000000_0111100101111000_0011110000000000"; -- 0.4744908809661865
	pesos_i(8915) := b"0000000000000000_0000000000000000_0100110011110111_1100011110000000"; -- 0.3006558120250702
	pesos_i(8916) := b"0000000000000000_0000000000000000_0011001010001000_1110101110000000"; -- 0.1974017322063446
	pesos_i(8917) := b"1111111111111111_1111111111111111_1100011011111101_1111001001000000"; -- -0.22268758714199066
	pesos_i(8918) := b"1111111111111111_1111111111111111_1011001100100101_1011100110000000"; -- -0.30020561814308167
	pesos_i(8919) := b"0000000000000000_0000000000000000_0000011000101001_0101000000110000"; -- 0.024067889899015427
	pesos_i(8920) := b"1111111111111111_1111111111111111_1001110000100011_1000101000000000"; -- -0.3900827169418335
	pesos_i(8921) := b"1111111111111111_1111111111111111_0111110011111000_0100011100000000"; -- -0.511836588382721
	pesos_i(8922) := b"0000000000000000_0000000000000000_0100011111100010_0100001010000000"; -- 0.28079620003700256
	pesos_i(8923) := b"1111111111111111_1111111111111111_1111011010101100_0010001110110000"; -- -0.03643586114048958
	pesos_i(8924) := b"0000000000000000_0000000000000000_1000100000100110_1111101100000000"; -- 0.5318447947502136
	pesos_i(8925) := b"1111111111111111_1111111111111111_0101100101110101_0110010100000000"; -- -0.6505524516105652
	pesos_i(8926) := b"1111111111111111_1111111111111110_1111011110101111_1111011000000000"; -- -1.0324712991714478
	pesos_i(8927) := b"0000000000000000_0000000000000000_1000010110010001_0111110000000000"; -- 0.5217511653900146
	pesos_i(8928) := b"1111111111111111_1111111111111111_1010110110010111_0001100100000000"; -- -0.3219131827354431
	pesos_i(8929) := b"0000000000000000_0000000000000000_0111101100001101_0110010000000000"; -- 0.48067307472229004
	pesos_i(8930) := b"1111111111111111_1111111111111111_1011111000100010_1011101010000000"; -- -0.2572825849056244
	pesos_i(8931) := b"1111111111111111_1111111111111111_1100010101001010_0101111010000000"; -- -0.22933396697044373
	pesos_i(8932) := b"0000000000000000_0000000000000000_0001011000011010_1110111111000000"; -- 0.0863485187292099
	pesos_i(8933) := b"0000000000000000_0000000000000000_0011101101100111_1111100011000000"; -- 0.23205523192882538
	pesos_i(8934) := b"1111111111111111_1111111111111111_1010000111101001_0010001000000000"; -- -0.36753642559051514
	pesos_i(8935) := b"1111111111111111_1111111111111111_1011101000000001_0010101110000000"; -- -0.27341964840888977
	pesos_i(8936) := b"0000000000000000_0000000000000000_0101010101101001_1100000110000000"; -- 0.33364495635032654
	pesos_i(8937) := b"1111111111111111_1111111111111111_1111011000000010_1011110100000000"; -- -0.03902071714401245
	pesos_i(8938) := b"0000000000000000_0000000000000000_0100111110000000_0100001110000000"; -- 0.31055089831352234
	pesos_i(8939) := b"0000000000000000_0000000000000000_0001110010110011_1001100110000000"; -- 0.11211547255516052
	pesos_i(8940) := b"1111111111111111_1111111111111111_0110000101011100_0101101000000000"; -- -0.6196845769882202
	pesos_i(8941) := b"0000000000000000_0000000000000000_0100011011010110_1110000100000000"; -- 0.27671629190444946
	pesos_i(8942) := b"1111111111111111_1111111111111111_1010100101010110_1000011010000000"; -- -0.3385234773159027
	pesos_i(8943) := b"0000000000000000_0000000000000000_0101000110000100_0011011110000000"; -- 0.31842371821403503
	pesos_i(8944) := b"1111111111111111_1111111111111111_1101100110000010_1111010010000000"; -- -0.15034553408622742
	pesos_i(8945) := b"0000000000000000_0000000000000000_0011101011110100_1110010101000000"; -- 0.23029930889606476
	pesos_i(8946) := b"0000000000000000_0000000000000000_0011000001110110_0100010010000000"; -- 0.18930462002754211
	pesos_i(8947) := b"1111111111111111_1111111111111111_1110101111000110_0110100100100000"; -- -0.07900374382734299
	pesos_i(8948) := b"0000000000000000_0000000000000000_0110010101100011_1111010110000000"; -- 0.39605650305747986
	pesos_i(8949) := b"0000000000000000_0000000000000000_0011001010001111_1110101010000000"; -- 0.19750848412513733
	pesos_i(8950) := b"0000000000000000_0000000000000000_0000011000000110_1111100110000000"; -- 0.02354392409324646
	pesos_i(8951) := b"1111111111111111_1111111111111110_1111100000000000_1001100000000000"; -- -1.0312409400939941
	pesos_i(8952) := b"1111111111111111_1111111111111111_1111100110000001_1001000001110000"; -- -0.025366757065057755
	pesos_i(8953) := b"0000000000000000_0000000000000000_0001010001101110_1100110101100000"; -- 0.07981570810079575
	pesos_i(8954) := b"0000000000000000_0000000000000000_0000111000110111_0001010010000000"; -- 0.055527955293655396
	pesos_i(8955) := b"1111111111111111_1111111111111111_1100100100011101_1000100110000000"; -- -0.21439304947853088
	pesos_i(8956) := b"1111111111111111_1111111111111111_1010010100101010_0000100110000000"; -- -0.35482731461524963
	pesos_i(8957) := b"1111111111111111_1111111111111111_1111011001011111_0010101000000000"; -- -0.037610411643981934
	pesos_i(8958) := b"1111111111111111_1111111111111111_1010111110111100_1010110110000000"; -- -0.31352725625038147
	pesos_i(8959) := b"1111111111111111_1111111111111111_1001011111111110_1011011000000000"; -- -0.4062696695327759
	pesos_i(8960) := b"0000000000000000_0000000000000000_0101001100101010_0011110010000000"; -- 0.3248632252216339
	pesos_i(8961) := b"1111111111111111_1111111111111111_1111100011000001_0001100000100000"; -- -0.028303615748882294
	pesos_i(8962) := b"0000000000000000_0000000000000000_0010000110101101_1011110101000000"; -- 0.13155730068683624
	pesos_i(8963) := b"1111111111111111_1111111111111111_0101101100000011_1111101000000000"; -- -0.6444705724716187
	pesos_i(8964) := b"0000000000000000_0000000000000000_0001010000101011_1111011101000000"; -- 0.07879586517810822
	pesos_i(8965) := b"0000000000000000_0000000000000000_0011111010000110_0000010110000000"; -- 0.24423250555992126
	pesos_i(8966) := b"1111111111111111_1111111111111111_1111110011000101_0010111001001000"; -- -0.012616259977221489
	pesos_i(8967) := b"1111111111111111_1111111111111111_1011110010000101_0000110110000000"; -- -0.26359477639198303
	pesos_i(8968) := b"1111111111111111_1111111111111111_1100100101101110_1000111010000000"; -- -0.2131567895412445
	pesos_i(8969) := b"0000000000000000_0000000000000000_0001010000101001_1101111001100000"; -- 0.07876386493444443
	pesos_i(8970) := b"0000000000000000_0000000000000000_0000110011110111_0001000001010000"; -- 0.0506448931992054
	pesos_i(8971) := b"0000000000000000_0000000000000000_0011110011101101_1010001111000000"; -- 0.23800109326839447
	pesos_i(8972) := b"1111111111111111_1111111111111110_1011000101001000_1111011000000000"; -- -1.3074804544448853
	pesos_i(8973) := b"0000000000000000_0000000000000001_0001111011010110_0011001000000000"; -- 1.1204558610916138
	pesos_i(8974) := b"1111111111111111_1111111111111111_1011001010101000_1010110100000000"; -- -0.30211371183395386
	pesos_i(8975) := b"1111111111111111_1111111111111111_1000111110110011_1101001100000000"; -- -0.4386623501777649
	pesos_i(8976) := b"0000000000000000_0000000000000000_0101100010011000_0100011000000000"; -- 0.3460735082626343
	pesos_i(8977) := b"0000000000000000_0000000000000000_0000000011111101_1111101011110001"; -- 0.0038754309061914682
	pesos_i(8978) := b"1111111111111111_1111111111111111_0110010101101011_0000000000000000"; -- -0.6038360595703125
	pesos_i(8979) := b"1111111111111111_1111111111111111_0111010001100101_0100000100000000"; -- -0.5453299880027771
	pesos_i(8980) := b"1111111111111111_1111111111111111_1110110110001001_1100010100000000"; -- -0.07211655378341675
	pesos_i(8981) := b"1111111111111111_1111111111111111_1111110101010101_1000011111111000"; -- -0.010413648560643196
	pesos_i(8982) := b"1111111111111111_1111111111111111_1110100001000010_0011010111000000"; -- -0.09273971617221832
	pesos_i(8983) := b"0000000000000000_0000000000000000_1000011111000000_0001111000000000"; -- 0.5302752256393433
	pesos_i(8984) := b"1111111111111111_1111111111111110_1010010111111001_1101011000000000"; -- -1.3516565561294556
	pesos_i(8985) := b"1111111111111111_1111111111111111_0111100001001101_0100110000000000"; -- -0.5300705432891846
	pesos_i(8986) := b"0000000000000000_0000000000000000_0010011010111001_1110101111000000"; -- 0.1512744277715683
	pesos_i(8987) := b"0000000000000000_0000000000000000_0000010100101011_1010111011000000"; -- 0.020197793841362
	pesos_i(8988) := b"0000000000000000_0000000000000000_0100001101010001_1011000110000000"; -- 0.26296529173851013
	pesos_i(8989) := b"1111111111111111_1111111111111111_0111010011100000_1010111100000000"; -- -0.5434466004371643
	pesos_i(8990) := b"1111111111111111_1111111111111111_1110110010111011_0011100110000000"; -- -0.07526817917823792
	pesos_i(8991) := b"0000000000000000_0000000000000000_0100111011010111_1011100110000000"; -- 0.30797919631004333
	pesos_i(8992) := b"1111111111111111_1111111111111111_1101001110010001_0011011010000000"; -- -0.17356547713279724
	pesos_i(8993) := b"1111111111111111_1111111111111111_0110100100110010_0111110000000000"; -- -0.5890734195709229
	pesos_i(8994) := b"0000000000000000_0000000000000000_0100010000001110_0001011010000000"; -- 0.26583996415138245
	pesos_i(8995) := b"1111111111111111_1111111111111111_1100110110110111_0110100110000000"; -- -0.1964201033115387
	pesos_i(8996) := b"0000000000000000_0000000000000000_0110100000010101_1101100010000000"; -- 0.40658333897590637
	pesos_i(8997) := b"1111111111111111_1111111111111111_0111010001111110_0001111000000000"; -- -0.5449506044387817
	pesos_i(8998) := b"1111111111111111_1111111111111111_1101101110000000_0010110101000000"; -- -0.1425754278898239
	pesos_i(8999) := b"0000000000000000_0000000000000000_0100100110001001_1111000110000000"; -- 0.28726109862327576
	pesos_i(9000) := b"1111111111111111_1111111111111111_1000011000010111_1000000110000000"; -- -0.4762038290500641
	pesos_i(9001) := b"0000000000000000_0000000000000000_0101011100111110_0111010100000000"; -- 0.3407967686653137
	pesos_i(9002) := b"1111111111111111_1111111111111111_0010011100000001_1111101100000000"; -- -0.8476260304450989
	pesos_i(9003) := b"0000000000000000_0000000000000000_0101000010111100_0101111110000000"; -- 0.31537434458732605
	pesos_i(9004) := b"1111111111111111_1111111111111111_1101010001110110_0101110110000000"; -- -0.1700688898563385
	pesos_i(9005) := b"0000000000000000_0000000000000000_0001011011001011_1000000010100000"; -- 0.08904270082712173
	pesos_i(9006) := b"1111111111111111_1111111111111111_0100000111011101_1011010000000000"; -- -0.7427108287811279
	pesos_i(9007) := b"0000000000000000_0000000000000000_1010100100000010_1011011000000000"; -- 0.6601976156234741
	pesos_i(9008) := b"1111111111111111_1111111111111111_1101110010100110_1100010111000000"; -- -0.13808025419712067
	pesos_i(9009) := b"1111111111111111_1111111111111111_1101111101000100_1101100011000000"; -- -0.12785573303699493
	pesos_i(9010) := b"1111111111111111_1111111111111111_0110011000011110_0011101000000000"; -- -0.601101279258728
	pesos_i(9011) := b"0000000000000000_0000000000000000_1001101110011100_1110010000000000"; -- 0.6078627109527588
	pesos_i(9012) := b"1111111111111111_1111111111111111_1100000111011011_1000001001000000"; -- -0.2427443116903305
	pesos_i(9013) := b"0000000000000000_0000000000000000_0001110000011111_1010111010100000"; -- 0.1098584309220314
	pesos_i(9014) := b"0000000000000000_0000000000000000_0001011101011010_1001010011100000"; -- 0.09122591465711594
	pesos_i(9015) := b"1111111111111111_1111111111111111_1011100110111100_1001000000000000"; -- -0.27446651458740234
	pesos_i(9016) := b"0000000000000000_0000000000000000_0100111011011111_1110100100000000"; -- 0.30810409784317017
	pesos_i(9017) := b"1111111111111111_1111111111111111_1100111100000001_1001100001000000"; -- -0.19138191640377045
	pesos_i(9018) := b"0000000000000000_0000000000000000_0101010001011011_0111101110000000"; -- 0.32952091097831726
	pesos_i(9019) := b"1111111111111111_1111111111111111_1000001010111000_0100111010000000"; -- -0.48937520384788513
	pesos_i(9020) := b"0000000000000000_0000000000000000_0000010011011101_0011010001011000"; -- 0.019000312313437462
	pesos_i(9021) := b"1111111111111111_1111111111111111_1000111101000010_1010101010000000"; -- -0.4403890073299408
	pesos_i(9022) := b"0000000000000000_0000000000000000_0010110000110111_1000101001000000"; -- 0.1727224737405777
	pesos_i(9023) := b"1111111111111111_1111111111111111_1000000010000001_1001001010000000"; -- -0.4980228841304779
	pesos_i(9024) := b"0000000000000000_0000000000000000_0011110001100011_0100000101000000"; -- 0.2358895093202591
	pesos_i(9025) := b"1111111111111111_1111111111111111_1000100111101011_1110010110000000"; -- -0.46124425530433655
	pesos_i(9026) := b"0000000000000000_0000000000000000_0101010111011110_0000001100000000"; -- 0.3354188799858093
	pesos_i(9027) := b"0000000000000000_0000000000000000_0010001010011111_1001001011000000"; -- 0.1352473944425583
	pesos_i(9028) := b"0000000000000000_0000000000000000_0110100100001101_1000011000000000"; -- 0.4103626012802124
	pesos_i(9029) := b"1111111111111111_1111111111111111_0011111101100111_0001000100000000"; -- -0.7523335814476013
	pesos_i(9030) := b"1111111111111111_1111111111111111_1111010001111111_1010010010100000"; -- -0.04492732137441635
	pesos_i(9031) := b"1111111111111111_1111111111111111_1100100100110001_1000010100000000"; -- -0.21408814191818237
	pesos_i(9032) := b"1111111111111111_1111111111111111_0011101001111110_0110100000000000"; -- -0.7715086936950684
	pesos_i(9033) := b"1111111111111111_1111111111111111_1100100011111010_0011110100000000"; -- -0.2149316668510437
	pesos_i(9034) := b"0000000000000000_0000000000000000_0000110000001101_0000000000110000"; -- 0.047073375433683395
	pesos_i(9035) := b"0000000000000000_0000000000000000_0000111111100101_0111010110100000"; -- 0.062095023691654205
	pesos_i(9036) := b"0000000000000000_0000000000000000_0101111011100000_0100100000000000"; -- 0.37060976028442383
	pesos_i(9037) := b"0000000000000000_0000000000000000_0000100111111011_1100010001000000"; -- 0.03899790346622467
	pesos_i(9038) := b"1111111111111111_1111111111111111_0111101101101111_1101000000000000"; -- -0.5178251266479492
	pesos_i(9039) := b"0000000000000000_0000000000000000_0011010101100001_1100101010000000"; -- 0.20852342247962952
	pesos_i(9040) := b"0000000000000000_0000000000000000_0010110011010010_1111110011000000"; -- 0.17509441077709198
	pesos_i(9041) := b"1111111111111111_1111111111111111_1011011011001111_1110001110000000"; -- -0.2858903706073761
	pesos_i(9042) := b"0000000000000000_0000000000000000_0000010101101101_1100101011000000"; -- 0.02120654284954071
	pesos_i(9043) := b"1111111111111111_1111111111111111_1010000101001111_0110111000000000"; -- -0.3698817491531372
	pesos_i(9044) := b"1111111111111111_1111111111111111_1011000111111111_0000010100000000"; -- -0.3047024607658386
	pesos_i(9045) := b"0000000000000000_0000000000000000_0011001001100000_0000110010000000"; -- 0.1967780888080597
	pesos_i(9046) := b"0000000000000000_0000000000000000_0100011100101010_1001101110000000"; -- 0.2779938876628876
	pesos_i(9047) := b"0000000000000000_0000000000000000_0011111110110101_0111001101000000"; -- 0.24886246025562286
	pesos_i(9048) := b"1111111111111111_1111111111111111_1000101001110101_1010010010000000"; -- -0.45914241671562195
	pesos_i(9049) := b"0000000000000000_0000000000000000_0011011100000111_0010100111000000"; -- 0.21495305001735687
	pesos_i(9050) := b"0000000000000000_0000000000000000_0010100101011010_0001000110000000"; -- 0.16153058409690857
	pesos_i(9051) := b"1111111111111111_1111111111111111_1111101101111001_0111011000101000"; -- -0.017677893862128258
	pesos_i(9052) := b"0000000000000000_0000000000000000_0111111011011000_0101100110000000"; -- 0.4954887330532074
	pesos_i(9053) := b"1111111111111111_1111111111111111_0110110001100100_0100000100000000"; -- -0.5765952467918396
	pesos_i(9054) := b"1111111111111111_1111111111111111_1110010111111000_0110000000000000"; -- -0.10167884826660156
	pesos_i(9055) := b"0000000000000000_0000000000000000_0000010011000000_1111001110100000"; -- 0.018569208681583405
	pesos_i(9056) := b"0000000000000000_0000000000000000_0101011010000100_1011111000000000"; -- 0.3379629850387573
	pesos_i(9057) := b"1111111111111111_1111111111111111_1100101101100010_1010010001000000"; -- -0.20552609860897064
	pesos_i(9058) := b"1111111111111111_1111111111111111_1010101100100000_0101010100000000"; -- -0.3315379023551941
	pesos_i(9059) := b"0000000000000000_0000000000000000_0011010101101000_1100011110000000"; -- 0.2086300551891327
	pesos_i(9060) := b"1111111111111111_1111111111111111_1001000001111001_1011100100000000"; -- -0.43564265966415405
	pesos_i(9061) := b"0000000000000000_0000000000000000_0100100000111101_0001001000000000"; -- 0.28218185901641846
	pesos_i(9062) := b"1111111111111111_1111111111111111_0100001100000111_0111111100000000"; -- -0.738166868686676
	pesos_i(9063) := b"0000000000000000_0000000000000000_0001101110101010_0111000010000000"; -- 0.10806944966316223
	pesos_i(9064) := b"0000000000000000_0000000000000000_1100010111111000_1010111100000000"; -- 0.7733258605003357
	pesos_i(9065) := b"1111111111111111_1111111111111111_1001101001101000_0010100000000000"; -- -0.396848201751709
	pesos_i(9066) := b"1111111111111111_1111111111111111_1110000010011010_1010000010000000"; -- -0.12264057993888855
	pesos_i(9067) := b"1111111111111111_1111111111111111_1000110101011001_1011001010000000"; -- -0.4478500783443451
	pesos_i(9068) := b"1111111111111111_1111111111111111_1111001111011010_1110010001100000"; -- -0.04744122177362442
	pesos_i(9069) := b"0000000000000000_0000000000000000_1010011110000010_1001010100000000"; -- 0.6543362736701965
	pesos_i(9070) := b"1111111111111111_1111111111111111_0100001110010001_1100101000000000"; -- -0.7360566854476929
	pesos_i(9071) := b"1111111111111111_1111111111111111_0101011001101000_1101110100000000"; -- -0.6624624133110046
	pesos_i(9072) := b"0000000000000000_0000000000000000_0111000110010101_1101000100000000"; -- 0.44369226694107056
	pesos_i(9073) := b"1111111111111111_1111111111111111_1000011101010011_0100100110000000"; -- -0.4713853895664215
	pesos_i(9074) := b"1111111111111111_1111111111111111_1010110100100111_0011010110000000"; -- -0.323620468378067
	pesos_i(9075) := b"0000000000000000_0000000000000000_0011010001010001_0110010011000000"; -- 0.20436696708202362
	pesos_i(9076) := b"1111111111111111_1111111111111111_0111110110001011_0110101000000000"; -- -0.5095914602279663
	pesos_i(9077) := b"0000000000000000_0000000000000000_0010011000010100_0000110110000000"; -- 0.14874348044395447
	pesos_i(9078) := b"1111111111111111_1111111111111111_0110000100010110_1110000100000000"; -- -0.6207446455955505
	pesos_i(9079) := b"0000000000000000_0000000000000000_0001101100100010_0010010110100000"; -- 0.10598979145288467
	pesos_i(9080) := b"1111111111111111_1111111111111111_1010111000101001_0111110000000000"; -- -0.31967949867248535
	pesos_i(9081) := b"0000000000000000_0000000000000000_0010001010101000_1101111010000000"; -- 0.13538923859596252
	pesos_i(9082) := b"0000000000000000_0000000000000000_0011101101110111_0100010101000000"; -- 0.2322886735200882
	pesos_i(9083) := b"1111111111111111_1111111111111111_0111000000011111_0110000000000000"; -- -0.5620212554931641
	pesos_i(9084) := b"1111111111111111_1111111111111111_1101000110011111_1011111111000000"; -- -0.18115617334842682
	pesos_i(9085) := b"0000000000000000_0000000000000000_0010111100100010_0000001101000000"; -- 0.18411274254322052
	pesos_i(9086) := b"0000000000000000_0000000000000000_0001101100010001_1101011110000000"; -- 0.1057409942150116
	pesos_i(9087) := b"1111111111111111_1111111111111111_1110100011101110_1111100111100000"; -- -0.09010351449251175
	pesos_i(9088) := b"0000000000000000_0000000000000000_0000101001000001_1101000101110000"; -- 0.040066804736852646
	pesos_i(9089) := b"1111111111111111_1111111111111111_1010101111100111_1011110000000000"; -- -0.3284952640533447
	pesos_i(9090) := b"1111111111111111_1111111111111111_1110001110110000_0100000010100000"; -- -0.11059185117483139
	pesos_i(9091) := b"1111111111111111_1111111111111111_1010011010000000_0100000010000000"; -- -0.349605530500412
	pesos_i(9092) := b"0000000000000000_0000000000000000_0010010010110110_1101010001000000"; -- 0.14341475069522858
	pesos_i(9093) := b"1111111111111111_1111111111111111_1100100100111001_0101100101000000"; -- -0.2139686793088913
	pesos_i(9094) := b"1111111111111111_1111111111111111_1111100011101101_0100001111101000"; -- -0.02762961946427822
	pesos_i(9095) := b"1111111111111111_1111111111111111_1111100001001111_1111111001100000"; -- -0.03002939373254776
	pesos_i(9096) := b"0000000000000000_0000000000000000_0100000010010111_1111001010000000"; -- 0.25231853127479553
	pesos_i(9097) := b"1111111111111111_1111111111111111_0011101101110000_1011101000000000"; -- -0.7678111791610718
	pesos_i(9098) := b"1111111111111111_1111111111111111_1010101001001101_1001010010000000"; -- -0.33475372195243835
	pesos_i(9099) := b"1111111111111111_1111111111111111_1101010101010001_1000110000000000"; -- -0.16672444343566895
	pesos_i(9100) := b"0000000000000000_0000000000000000_0010101001011110_0100111101000000"; -- 0.16550154983997345
	pesos_i(9101) := b"0000000000000000_0000000000000000_0011110001100000_0001101001000000"; -- 0.23584140837192535
	pesos_i(9102) := b"0000000000000000_0000000000000000_0000100001110101_1110000000110000"; -- 0.03304864093661308
	pesos_i(9103) := b"1111111111111111_1111111111111111_1111101010100011_1100000110011000"; -- -0.020938778296113014
	pesos_i(9104) := b"0000000000000000_0000000000000000_0101100001111100_1010001010000000"; -- 0.345651775598526
	pesos_i(9105) := b"1111111111111111_1111111111111111_1101111110011111_0000001100000000"; -- -0.12647992372512817
	pesos_i(9106) := b"1111111111111111_1111111111111111_1110011101010101_0110100001100000"; -- -0.09635303169488907
	pesos_i(9107) := b"1111111111111111_1111111111111111_1111100000111111_1101010001101000"; -- -0.030276035889983177
	pesos_i(9108) := b"1111111111111111_1111111111111111_1000000100000101_1011011000000000"; -- -0.4960066080093384
	pesos_i(9109) := b"0000000000000000_0000000000000000_1000000111011011_0000011000000000"; -- 0.5072482824325562
	pesos_i(9110) := b"1111111111111111_1111111111111111_1011100100101110_1001100110000000"; -- -0.276632696390152
	pesos_i(9111) := b"0000000000000000_0000000000000000_0011101110110111_0101010100000000"; -- 0.2332661747932434
	pesos_i(9112) := b"1111111111111111_1111111111111111_1001101001110010_1011010110000000"; -- -0.39668717980384827
	pesos_i(9113) := b"0000000000000000_0000000000000000_0001011011001000_0010001110100000"; -- 0.08899138122797012
	pesos_i(9114) := b"0000000000000000_0000000000000000_0101011100101110_0010011110000000"; -- 0.34054800868034363
	pesos_i(9115) := b"1111111111111111_1111111111111111_0001000011110110_0011000000000000"; -- -0.9337434768676758
	pesos_i(9116) := b"0000000000000000_0000000000000000_0000000100111110_1000101110100010"; -- 0.004860617686063051
	pesos_i(9117) := b"1111111111111111_1111111111111111_1010101011001110_0011101100000000"; -- -0.33279067277908325
	pesos_i(9118) := b"0000000000000000_0000000000000000_0010110111011110_0010011011000000"; -- 0.17917101085186005
	pesos_i(9119) := b"0000000000000000_0000000000000000_1110010010100100_0001101000000000"; -- 0.8931289911270142
	pesos_i(9120) := b"1111111111111111_1111111111111111_0101000101100110_1110100100000000"; -- -0.6820234656333923
	pesos_i(9121) := b"1111111111111111_1111111111111111_1001011000010110_1010100110000000"; -- -0.41371670365333557
	pesos_i(9122) := b"1111111111111111_1111111111111111_1011100100100100_1110000000000000"; -- -0.2767810821533203
	pesos_i(9123) := b"1111111111111111_1111111111111111_1000011100010100_1111111110000000"; -- -0.4723358452320099
	pesos_i(9124) := b"0000000000000000_0000000000000000_0000110111011100_0100100111100000"; -- 0.05414258688688278
	pesos_i(9125) := b"1111111111111111_1111111111111111_1010110110011110_0101000010000000"; -- -0.3218030631542206
	pesos_i(9126) := b"0000000000000000_0000000000000000_0010111111000011_1100101000000000"; -- 0.18658125400543213
	pesos_i(9127) := b"1111111111111111_1111111111111111_1100111001111101_0110110101000000"; -- -0.1933986395597458
	pesos_i(9128) := b"1111111111111111_1111111111111111_1010101111100100_0100110010000000"; -- -0.3285476863384247
	pesos_i(9129) := b"1111111111111111_1111111111111111_1111010111100010_0111100101100000"; -- -0.03951302915811539
	pesos_i(9130) := b"0000000000000000_0000000000000000_0011100001110010_0011010101000000"; -- 0.2204926759004593
	pesos_i(9131) := b"0000000000000000_0000000000000000_0010111010001010_0110101110000000"; -- 0.18179962038993835
	pesos_i(9132) := b"1111111111111111_1111111111111111_1010011100011010_1110110110000000"; -- -0.34724536538124084
	pesos_i(9133) := b"1111111111111111_1111111111111111_1011100111011101_1010001110000000"; -- -0.2739618122577667
	pesos_i(9134) := b"1111111111111111_1111111111111111_1001001001001010_0011010110000000"; -- -0.4285551607608795
	pesos_i(9135) := b"0000000000000000_0000000000000000_0001101101110110_0101100100000000"; -- 0.10727459192276001
	pesos_i(9136) := b"1111111111111111_1111111111111111_1100111101110010_1001110100000000"; -- -0.18965739011764526
	pesos_i(9137) := b"1111111111111111_1111111111111111_1011100000101101_0010011110000000"; -- -0.28056100010871887
	pesos_i(9138) := b"0000000000000000_0000000000000000_0100010000101000_1001111100000000"; -- 0.2662448287010193
	pesos_i(9139) := b"1111111111111111_1111111111111111_1101111001100111_0111011000000000"; -- -0.131233811378479
	pesos_i(9140) := b"0000000000000000_0000000000000000_0010111010111110_1011010100000000"; -- 0.18259745836257935
	pesos_i(9141) := b"0000000000000000_0000000000000000_0010011010100110_1101110101000000"; -- 0.15098364651203156
	pesos_i(9142) := b"1111111111111111_1111111111111111_1111111101110111_1000110110010010"; -- -0.0020820158533751965
	pesos_i(9143) := b"0000000000000000_0000000000000000_0010011011000010_0010001001000000"; -- 0.15139974653720856
	pesos_i(9144) := b"0000000000000000_0000000000000000_0011010010110101_1010101111000000"; -- 0.20589707791805267
	pesos_i(9145) := b"0000000000000000_0000000000000000_0000011000010101_0101100001100000"; -- 0.023763202130794525
	pesos_i(9146) := b"1111111111111111_1111111111111111_1110101110001011_0000110111100000"; -- -0.07990945130586624
	pesos_i(9147) := b"1111111111111111_1111111111111111_1000000010111001_1111011110000000"; -- -0.4971623718738556
	pesos_i(9148) := b"1111111111111111_1111111111111111_1111000100100111_0101010110010000"; -- -0.057993557304143906
	pesos_i(9149) := b"1111111111111111_1111111111111111_1001000001000001_1001111010000000"; -- -0.4364987313747406
	pesos_i(9150) := b"1111111111111111_1111111111111111_1001101111000110_0101100100000000"; -- -0.39150470495224
	pesos_i(9151) := b"0000000000000000_0000000000000000_0000000010011000_1001001000111000"; -- 0.0023280512541532516
	pesos_i(9152) := b"1111111111111111_1111111111111111_0110111011011111_1111100000000000"; -- -0.5668950080871582
	pesos_i(9153) := b"0000000000000000_0000000000000000_0101111110000001_1000011000000000"; -- 0.3730701208114624
	pesos_i(9154) := b"0000000000000000_0000000000000000_0101100101101100_1010101110000000"; -- 0.349314421415329
	pesos_i(9155) := b"0000000000000000_0000000000000000_0000011101110111_0111101110001000"; -- 0.02916690893471241
	pesos_i(9156) := b"1111111111111111_1111111111111111_0111110010111101_1010001000000000"; -- -0.5127314329147339
	pesos_i(9157) := b"0000000000000000_0000000000000000_0001101101000111_1101000011000000"; -- 0.10656456649303436
	pesos_i(9158) := b"1111111111111111_1111111111111111_0111011100111111_0110001100000000"; -- -0.5341890454292297
	pesos_i(9159) := b"1111111111111111_1111111111111111_1110110100010100_1011001001000000"; -- -0.07390294969081879
	pesos_i(9160) := b"0000000000000000_0000000000000000_0010110101110010_0111111000000000"; -- 0.1775282621383667
	pesos_i(9161) := b"0000000000000000_0000000000000000_0000010010011001_0000001001001000"; -- 0.017959730699658394
	pesos_i(9162) := b"0000000000000000_0000000000000000_0001001110100111_1110100100100000"; -- 0.07678086310625076
	pesos_i(9163) := b"1111111111111111_1111111111111111_1111101001100101_1101111000101000"; -- -0.021883120760321617
	pesos_i(9164) := b"0000000000000000_0000000000000000_0000110100001000_1011101101100000"; -- 0.05091448873281479
	pesos_i(9165) := b"1111111111111111_1111111111111111_1101101011010110_1111100110000000"; -- -0.14515724778175354
	pesos_i(9166) := b"0000000000000000_0000000000000000_0001010010110010_0100010010000000"; -- 0.08084514737129211
	pesos_i(9167) := b"0000000000000000_0000000000000000_0000001110001001_0001000010010100"; -- 0.013810192234814167
	pesos_i(9168) := b"0000000000000000_0000000000000000_0010010111001001_1100000111000000"; -- 0.14760981500148773
	pesos_i(9169) := b"1111111111111111_1111111111111111_1101110110110111_0011111001000000"; -- -0.13392268121242523
	pesos_i(9170) := b"0000000000000000_0000000000000000_0000011001001110_1011101110001000"; -- 0.024638863280415535
	pesos_i(9171) := b"0000000000000000_0000000000000000_0000001011000000_1000011110010100"; -- 0.010750268585979939
	pesos_i(9172) := b"0000000000000000_0000000000000000_0000010100000101_0101001101010000"; -- 0.01961250975728035
	pesos_i(9173) := b"1111111111111111_1111111111111111_0011111111001000_1110000100000000"; -- -0.7508410811424255
	pesos_i(9174) := b"1111111111111111_1111111111111111_1110000110101110_0001110101100000"; -- -0.11843696981668472
	pesos_i(9175) := b"0000000000000000_0000000000000000_0011111100101011_0001110110000000"; -- 0.24675163626670837
	pesos_i(9176) := b"1111111111111111_1111111111111111_1001000110110001_1001000010000000"; -- -0.43088433146476746
	pesos_i(9177) := b"1111111111111111_1111111111111111_1100010010111111_0001010111000000"; -- -0.23145927488803864
	pesos_i(9178) := b"1111111111111111_1111111111111111_1001110100100000_1111111100000000"; -- -0.3862152695655823
	pesos_i(9179) := b"0000000000000000_0000000000000000_0101010110111110_1110100100000000"; -- 0.33494430780410767
	pesos_i(9180) := b"0000000000000000_0000000000000000_0000011101000010_1111110111101000"; -- 0.0283659640699625
	pesos_i(9181) := b"0000000000000000_0000000000000000_0011011000100111_1101111001000000"; -- 0.21154583990573883
	pesos_i(9182) := b"1111111111111111_1111111111111111_0101101110111100_0001001000000000"; -- -0.641661524772644
	pesos_i(9183) := b"1111111111111111_1111111111111111_1100101110100101_0001111101000000"; -- -0.20451168715953827
	pesos_i(9184) := b"1111111111111111_1111111111111111_0011110100101100_0101000100000000"; -- -0.7610425353050232
	pesos_i(9185) := b"0000000000000000_0000000000000000_1000001011110011_0111001000000000"; -- 0.5115271806716919
	pesos_i(9186) := b"0000000000000000_0000000000000000_0010101010110111_1000011110000000"; -- 0.16686293482780457
	pesos_i(9187) := b"0000000000000000_0000000000000000_0110110100001001_0001000100000000"; -- 0.4259195923805237
	pesos_i(9188) := b"1111111111111111_1111111111111111_1100011111000110_0001101000000000"; -- -0.21963346004486084
	pesos_i(9189) := b"1111111111111111_1111111111111111_0001001111100100_0011110000000000"; -- -0.9222986698150635
	pesos_i(9190) := b"0000000000000000_0000000000000000_0000100011111010_1001010000100000"; -- 0.035073526203632355
	pesos_i(9191) := b"0000000000000000_0000000000000000_0101101000000101_0101101110000000"; -- 0.35164424777030945
	pesos_i(9192) := b"0000000000000000_0000000000000000_0100101011110010_1101101000000000"; -- 0.29276812076568604
	pesos_i(9193) := b"1111111111111111_1111111111111111_1011011000010000_0011000100000000"; -- -0.288815438747406
	pesos_i(9194) := b"1111111111111111_1111111111111111_1010111111010111_1101000010000000"; -- -0.31311318278312683
	pesos_i(9195) := b"0000000000000000_0000000000000000_0011110111100010_0111001110000000"; -- 0.24173662066459656
	pesos_i(9196) := b"1111111111111111_1111111111111111_1000100001010000_0101110000000000"; -- -0.46752381324768066
	pesos_i(9197) := b"1111111111111111_1111111111111111_1110001010000000_1101000101000000"; -- -0.11522190272808075
	pesos_i(9198) := b"1111111111111111_1111111111111111_0110001011100011_1110110100000000"; -- -0.6137096285820007
	pesos_i(9199) := b"1111111111111111_1111111111111111_1111101000100010_1111011011110000"; -- -0.022903982549905777
	pesos_i(9200) := b"0000000000000000_0000000000000000_0000111001001011_1010110111010000"; -- 0.05584226921200752
	pesos_i(9201) := b"0000000000000000_0000000000000000_0011001010111111_0010100000000000"; -- 0.19822931289672852
	pesos_i(9202) := b"0000000000000000_0000000000000000_1001111110101011_0111111100000000"; -- 0.623710572719574
	pesos_i(9203) := b"0000000000000000_0000000000000000_0000111100101100_1101000001000000"; -- 0.059277549386024475
	pesos_i(9204) := b"0000000000000000_0000000000000000_1001000110111111_0001000100000000"; -- 0.5693216919898987
	pesos_i(9205) := b"1111111111111111_1111111111111111_0010010000001000_1011100100000000"; -- -0.8592419028282166
	pesos_i(9206) := b"1111111111111111_1111111111111111_1101001101111110_1101100100000000"; -- -0.17384570837020874
	pesos_i(9207) := b"1111111111111111_1111111111111111_1110110100010100_1100111001100000"; -- -0.07390127331018448
	pesos_i(9208) := b"0000000000000000_0000000000000000_0101000011010000_0111010110000000"; -- 0.3156808316707611
	pesos_i(9209) := b"1111111111111111_1111111111111111_1001101000100010_0011101110000000"; -- -0.39791515469551086
	pesos_i(9210) := b"1111111111111111_1111111111111110_1101000010100100_1010011000000000"; -- -1.1849876642227173
	pesos_i(9211) := b"0000000000000000_0000000000000000_1000010010111111_0100111100000000"; -- 0.5185441374778748
	pesos_i(9212) := b"0000000000000000_0000000000000000_0000011010111001_0011100001000000"; -- 0.026263728737831116
	pesos_i(9213) := b"0000000000000000_0000000000000000_0100000110011001_1001001010000000"; -- 0.2562495768070221
	pesos_i(9214) := b"1111111111111111_1111111111111111_0111110011111111_1110010000000000"; -- -0.5117204189300537
	pesos_i(9215) := b"1111111111111111_1111111111111111_1101010011001000_1110100011000000"; -- -0.16880936920642853
	pesos_i(9216) := b"1111111111111111_1111111111111111_1111001010011101_0101100100100000"; -- -0.05228655785322189
	pesos_i(9217) := b"0000000000000000_0000000000000000_0110011000101101_1111110110000000"; -- 0.39913925528526306
	pesos_i(9218) := b"1111111111111111_1111111111111111_1011110100001100_0100000010000000"; -- -0.261531800031662
	pesos_i(9219) := b"1111111111111111_1111111111111111_1000011000100110_1101101110000000"; -- -0.4759695827960968
	pesos_i(9220) := b"0000000000000000_0000000000000000_0000010111011010_1111000011001000"; -- 0.022872017696499825
	pesos_i(9221) := b"1111111111111111_1111111111111111_1000010101001110_0111011010000000"; -- -0.4792715013027191
	pesos_i(9222) := b"1111111111111111_1111111111111111_0001111001111010_0010000000000000"; -- -0.8809490203857422
	pesos_i(9223) := b"0000000000000000_0000000000000000_0101011111101001_0110001110000000"; -- 0.34340497851371765
	pesos_i(9224) := b"0000000000000000_0000000000000000_1010001010111111_1011010000000000"; -- 0.6357376575469971
	pesos_i(9225) := b"0000000000000000_0000000000000000_0011110100001011_0011001110000000"; -- 0.23845216631889343
	pesos_i(9226) := b"1111111111111111_1111111111111111_1010110111010101_1011000010000000"; -- -0.32095810770988464
	pesos_i(9227) := b"1111111111111111_1111111111111111_0011001100101010_0111000000000000"; -- -0.8001337051391602
	pesos_i(9228) := b"1111111111111111_1111111111111111_0000010000101000_1111000100000000"; -- -0.9837502837181091
	pesos_i(9229) := b"0000000000000000_0000000000000000_1011001111010000_0011111100000000"; -- 0.7023963332176208
	pesos_i(9230) := b"1111111111111111_1111111111111111_0100101111001111_0010010000000000"; -- -0.7038705348968506
	pesos_i(9231) := b"1111111111111111_1111111111111111_0101010011110011_0101010100000000"; -- -0.6681620478630066
	pesos_i(9232) := b"1111111111111111_1111111111111111_1011011110111010_0000011100000000"; -- -0.2823176980018616
	pesos_i(9233) := b"1111111111111111_1111111111111111_0111100000101011_0110000000000000"; -- -0.5305881500244141
	pesos_i(9234) := b"1111111111111111_1111111111111111_1100100000011010_0010111000000000"; -- -0.21835052967071533
	pesos_i(9235) := b"1111111111111111_1111111111111111_1011111000011010_1001010010000000"; -- -0.25740692019462585
	pesos_i(9236) := b"0000000000000000_0000000000000000_0111111000111101_1011000100000000"; -- 0.49312883615493774
	pesos_i(9237) := b"0000000000000000_0000000000000000_0010001011010110_0011110101000000"; -- 0.1360815316438675
	pesos_i(9238) := b"1111111111111111_1111111111111111_1111101011010001_0000100011000000"; -- -0.020247891545295715
	pesos_i(9239) := b"1111111111111111_1111111111111111_1001000110001101_0101110010000000"; -- -0.4314367473125458
	pesos_i(9240) := b"0000000000000000_0000000000000000_0011001111000101_0010100111000000"; -- 0.20222721993923187
	pesos_i(9241) := b"0000000000000000_0000000000000000_0011010101011110_1101100000000000"; -- 0.20847845077514648
	pesos_i(9242) := b"1111111111111111_1111111111111111_0101111011010000_0001011000000000"; -- -0.6296373605728149
	pesos_i(9243) := b"0000000000000000_0000000000000000_1000110011000010_1001101000000000"; -- 0.5498443841934204
	pesos_i(9244) := b"1111111111111111_1111111111111111_0001110000000100_0100001100000000"; -- -0.89055997133255
	pesos_i(9245) := b"1111111111111111_1111111111111111_1000110100011111_0011111110000000"; -- -0.44874194264411926
	pesos_i(9246) := b"0000000000000000_0000000000000000_0010001001011001_1011100001000000"; -- 0.13418151438236237
	pesos_i(9247) := b"0000000000000000_0000000000000000_0111000101110100_0101111110000000"; -- 0.44318196177482605
	pesos_i(9248) := b"0000000000000000_0000000000000000_1001011010110000_1001011100000000"; -- 0.5886320471763611
	pesos_i(9249) := b"0000000000000000_0000000000000000_0110000011100100_0000101100000000"; -- 0.37847965955734253
	pesos_i(9250) := b"1111111111111111_1111111111111111_1001100101011000_1111001000000000"; -- -0.40098655223846436
	pesos_i(9251) := b"1111111111111111_1111111111111111_1011001100001111_0000101100000000"; -- -0.30055171251296997
	pesos_i(9252) := b"1111111111111111_1111111111111111_1100100001000110_0000111111000000"; -- -0.2176809459924698
	pesos_i(9253) := b"0000000000000000_0000000000000000_0101010101001100_1101100010000000"; -- 0.33320382237434387
	pesos_i(9254) := b"1111111111111111_1111111111111111_1010010110101111_0011001110000000"; -- -0.35279539227485657
	pesos_i(9255) := b"0000000000000000_0000000000000000_0101000100000001_0000001100000000"; -- 0.3164216876029968
	pesos_i(9256) := b"1111111111111111_1111111111111110_1110101111110100_1101110000000000"; -- -1.0782949924468994
	pesos_i(9257) := b"0000000000000000_0000000000000000_1111010111010011_1110110000000000"; -- 0.9602649211883545
	pesos_i(9258) := b"1111111111111111_1111111111111111_0101111010111111_0010010100000000"; -- -0.6298958659172058
	pesos_i(9259) := b"1111111111111111_1111111111111111_1101000011100000_1101111011000000"; -- -0.18406875431537628
	pesos_i(9260) := b"1111111111111111_1111111111111110_0110000010100010_1110100000000000"; -- -1.622514247894287
	pesos_i(9261) := b"0000000000000000_0000000000000000_0000101111010100_0011100000100000"; -- 0.04620695859193802
	pesos_i(9262) := b"0000000000000000_0000000000000000_0111010001101010_1100100000000000"; -- 0.4547543525695801
	pesos_i(9263) := b"1111111111111111_1111111111111111_0111010010111101_0110001100000000"; -- -0.5439851880073547
	pesos_i(9264) := b"0000000000000000_0000000000000000_0101000111000110_0001000110000000"; -- 0.31942853331565857
	pesos_i(9265) := b"1111111111111111_1111111111111111_1110110010001010_0111111001000000"; -- -0.0760117620229721
	pesos_i(9266) := b"1111111111111111_1111111111111111_1100111001110011_1101111011000000"; -- -0.19354446232318878
	pesos_i(9267) := b"1111111111111111_1111111111111111_1111001001110110_0001001000010000"; -- -0.052885886281728745
	pesos_i(9268) := b"1111111111111111_1111111111111111_1110101000011010_0111011001000000"; -- -0.08553372323513031
	pesos_i(9269) := b"1111111111111111_1111111111111111_0110111101001000_1100111100000000"; -- -0.5652952790260315
	pesos_i(9270) := b"1111111111111111_1111111111111111_1100111110010010_1001110110000000"; -- -0.18916907906532288
	pesos_i(9271) := b"1111111111111111_1111111111111111_1010101010000111_0110111000000000"; -- -0.3338710069656372
	pesos_i(9272) := b"1111111111111111_1111111111111110_1110100000011010_1001000000000000"; -- -1.0933446884155273
	pesos_i(9273) := b"1111111111111111_1111111111111111_1110010000010000_1011101110100000"; -- -0.10911967605352402
	pesos_i(9274) := b"0000000000000000_0000000000000000_0101011001011101_1010100010000000"; -- 0.33736661076545715
	pesos_i(9275) := b"0000000000000000_0000000000000000_0001010000110010_0111001000000000"; -- 0.0788947343826294
	pesos_i(9276) := b"0000000000000000_0000000000000000_0001110000110011_1010101100100000"; -- 0.11016339808702469
	pesos_i(9277) := b"0000000000000000_0000000000000000_0010001000001110_1011100010000000"; -- 0.13303712010383606
	pesos_i(9278) := b"0000000000000000_0000000000000000_1001000111100111_1011001100000000"; -- 0.5699416995048523
	pesos_i(9279) := b"0000000000000000_0000000000000000_0000010000001110_0010010101000000"; -- 0.015840843319892883
	pesos_i(9280) := b"1111111111111111_1111111111111111_0110001001110000_0001010000000000"; -- -0.6154773235321045
	pesos_i(9281) := b"1111111111111111_1111111111111110_1110010010010110_0000110000000000"; -- -1.1070854663848877
	pesos_i(9282) := b"0000000000000000_0000000000000000_0011001111100010_1000001010000000"; -- 0.2026750147342682
	pesos_i(9283) := b"1111111111111111_1111111111111111_0111111010011000_0000111100000000"; -- -0.5054922699928284
	pesos_i(9284) := b"1111111111111111_1111111111111111_1011110100010001_0101100010000000"; -- -0.2614540755748749
	pesos_i(9285) := b"1111111111111111_1111111111111111_1111011110101011_1110001010010000"; -- -0.032533492892980576
	pesos_i(9286) := b"0000000000000000_0000000000000000_0010101010111001_0100110110000000"; -- 0.1668899953365326
	pesos_i(9287) := b"0000000000000000_0000000000000000_0111101000001110_1110110100000000"; -- 0.47679024934768677
	pesos_i(9288) := b"0000000000000000_0000000000000000_0100010011100101_1010101010000000"; -- 0.2691294252872467
	pesos_i(9289) := b"1111111111111111_1111111111111111_1110110000100111_0100011111000000"; -- -0.07752563059329987
	pesos_i(9290) := b"1111111111111111_1111111111111111_1001100101000100_0100111000000000"; -- -0.4013015031814575
	pesos_i(9291) := b"0000000000000000_0000000000000000_0011011101111101_1010001111000000"; -- 0.21676085889339447
	pesos_i(9292) := b"0000000000000000_0000000000000000_0101001110010101_0000001100000000"; -- 0.3264924883842468
	pesos_i(9293) := b"0000000000000000_0000000000000000_0010111001100101_0101100101000000"; -- 0.1812339574098587
	pesos_i(9294) := b"0000000000000000_0000000000000000_0001100110000110_0001111011100000"; -- 0.09970276802778244
	pesos_i(9295) := b"1111111111111111_1111111111111111_1101110011011111_1100001111000000"; -- -0.13721062242984772
	pesos_i(9296) := b"1111111111111111_1111111111111111_1011101111010000_1110010100000000"; -- -0.26634377241134644
	pesos_i(9297) := b"1111111111111111_1111111111111111_0111101101111011_0010101100000000"; -- -0.5176518559455872
	pesos_i(9298) := b"0000000000000000_0000000000000000_0000000110111100_0111100001100100"; -- 0.006782078184187412
	pesos_i(9299) := b"0000000000000000_0000000000000000_0101001101011001_1011100110000000"; -- 0.32558783888816833
	pesos_i(9300) := b"1111111111111111_1111111111111111_1011001010011110_0000000110000000"; -- -0.30227652192115784
	pesos_i(9301) := b"0000000000000000_0000000000000000_0000001011000111_1101001001100100"; -- 0.010861539281904697
	pesos_i(9302) := b"0000000000000000_0000000000000000_0100100000101111_0100010000000000"; -- 0.2819712162017822
	pesos_i(9303) := b"0000000000000000_0000000000000000_0010010100101110_1111100111000000"; -- 0.14524804055690765
	pesos_i(9304) := b"0000000000000000_0000000000000000_1010111111110000_0111010000000000"; -- 0.687262773513794
	pesos_i(9305) := b"1111111111111111_1111111111111111_1100101101100100_1000011111000000"; -- -0.20549727976322174
	pesos_i(9306) := b"1111111111111111_1111111111111111_0011000000011000_0000000000000000"; -- -0.8121337890625
	pesos_i(9307) := b"1111111111111111_1111111111111111_1001101110100011_0010001110000000"; -- -0.392041951417923
	pesos_i(9308) := b"1111111111111111_1111111111111111_0110010110000110_1100000000000000"; -- -0.6034126281738281
	pesos_i(9309) := b"0000000000000000_0000000000000000_0111001001100100_0111011000000000"; -- 0.4468454122543335
	pesos_i(9310) := b"0000000000000000_0000000000000000_0011001001011010_1100001111000000"; -- 0.19669745862483978
	pesos_i(9311) := b"1111111111111111_1111111111111111_1011111000101011_1001000010000000"; -- -0.25714775919914246
	pesos_i(9312) := b"1111111111111111_1111111111111111_1010101011101010_0111100000000000"; -- -0.33235979080200195
	pesos_i(9313) := b"0000000000000000_0000000000000000_0111000111001111_1110111000000000"; -- 0.44457900524139404
	pesos_i(9314) := b"0000000000000000_0000000000000000_0010100101100101_1101100101000000"; -- 0.16171033680438995
	pesos_i(9315) := b"1111111111111111_1111111111111111_1010101110100110_0001100110000000"; -- -0.3294967710971832
	pesos_i(9316) := b"0000000000000000_0000000000000000_0011111000001010_1011100001000000"; -- 0.24235107004642487
	pesos_i(9317) := b"1111111111111111_1111111111111111_1110101110111110_1100011000000000"; -- -0.07912027835845947
	pesos_i(9318) := b"1111111111111111_1111111111111111_1110000011101000_1011000100100000"; -- -0.12144940346479416
	pesos_i(9319) := b"1111111111111111_1111111111111111_1011101011100001_0100000110000000"; -- -0.2700003683567047
	pesos_i(9320) := b"0000000000000000_0000000000000000_0011110001001100_1000000010000000"; -- 0.23554232716560364
	pesos_i(9321) := b"1111111111111111_1111111111111111_0010001111101101_0010001100000000"; -- -0.8596628308296204
	pesos_i(9322) := b"1111111111111111_1111111111111111_1001010011111100_0111000000000000"; -- -0.41802310943603516
	pesos_i(9323) := b"0000000000000000_0000000000000000_1010101011011100_0110001100000000"; -- 0.6674253344535828
	pesos_i(9324) := b"0000000000000000_0000000000000000_1000111011000101_1100010100000000"; -- 0.5577052235603333
	pesos_i(9325) := b"1111111111111111_1111111111111111_1110010000000001_0000010001000000"; -- -0.1093594878911972
	pesos_i(9326) := b"1111111111111111_1111111111111111_1010011010101110_1011111000000000"; -- -0.3488961458206177
	pesos_i(9327) := b"0000000000000000_0000000000000000_1001101100011100_1101011100000000"; -- 0.6059088110923767
	pesos_i(9328) := b"1111111111111111_1111111111111111_0010001101000111_0011001000000000"; -- -0.8621948957443237
	pesos_i(9329) := b"0000000000000000_0000000000000000_1100011000000010_0000000000000000"; -- 0.773468017578125
	pesos_i(9330) := b"1111111111111111_1111111111111111_0110100111001001_0100100100000000"; -- -0.5867723822593689
	pesos_i(9331) := b"1111111111111111_1111111111111111_0101011000000010_0011010100000000"; -- -0.6640288233757019
	pesos_i(9332) := b"1111111111111111_1111111111111111_0101111101000011_0001000100000000"; -- -0.6278828978538513
	pesos_i(9333) := b"1111111111111111_1111111111111111_0111011111011100_0010000100000000"; -- -0.5317973494529724
	pesos_i(9334) := b"0000000000000000_0000000000000000_0011110111011000_0100100101000000"; -- 0.2415815144777298
	pesos_i(9335) := b"1111111111111111_1111111111111111_1101110011011000_1010110111000000"; -- -0.13731874525547028
	pesos_i(9336) := b"0000000000000000_0000000000000000_0100011000000100_0111010000000000"; -- 0.27350544929504395
	pesos_i(9337) := b"0000000000000000_0000000000000000_0000101000101100_1100010010000000"; -- 0.039745599031448364
	pesos_i(9338) := b"0000000000000000_0000000000000000_0110000101000011_1000011010000000"; -- 0.3799366056919098
	pesos_i(9339) := b"0000000000000000_0000000000000000_0011111101001101_0011100111000000"; -- 0.24727211892604828
	pesos_i(9340) := b"1111111111111111_1111111111111111_1111101011010110_0111011101011000"; -- -0.020165005698800087
	pesos_i(9341) := b"1111111111111111_1111111111111111_0011011000010111_0000100000000000"; -- -0.7887110710144043
	pesos_i(9342) := b"1111111111111111_1111111111111111_1010100110110001_0110010000000000"; -- -0.33713698387145996
	pesos_i(9343) := b"1111111111111111_1111111111111111_1110111011011101_1000010101100000"; -- -0.06693235784769058
	pesos_i(9344) := b"0000000000000000_0000000000000000_0010101000011110_1100101110000000"; -- 0.1645323932170868
	pesos_i(9345) := b"0000000000000000_0000000000000000_0010011001000110_1011010101000000"; -- 0.14951641857624054
	pesos_i(9346) := b"0000000000000000_0000000000000000_0111001001000010_0001100010000000"; -- 0.446321040391922
	pesos_i(9347) := b"1111111111111111_1111111111111111_0110010110101100_1101110100000000"; -- -0.6028310656547546
	pesos_i(9348) := b"1111111111111111_1111111111111111_1010110000010010_0101011000000000"; -- -0.3278452157974243
	pesos_i(9349) := b"0000000000000000_0000000000000000_0110100111111000_0001001000000000"; -- 0.41394150257110596
	pesos_i(9350) := b"1111111111111111_1111111111111110_1111000100001101_1101111000000000"; -- -1.0583821535110474
	pesos_i(9351) := b"0000000000000000_0000000000000000_0011000011010010_1111011110000000"; -- 0.1907190978527069
	pesos_i(9352) := b"1111111111111111_1111111111111111_1010110000001100_1011010100000000"; -- -0.32793110609054565
	pesos_i(9353) := b"0000000000000000_0000000000000000_0011011010011111_1001011011000000"; -- 0.2133726328611374
	pesos_i(9354) := b"0000000000000000_0000000000000000_0000110111001010_0001110111000000"; -- 0.05386529862880707
	pesos_i(9355) := b"1111111111111111_1111111111111111_0111111001111011_1111111000000000"; -- -0.5059205293655396
	pesos_i(9356) := b"0000000000000000_0000000000000000_0011010100111010_1001101111000000"; -- 0.20792554318904877
	pesos_i(9357) := b"1111111111111111_1111111111111111_1110111001110001_1011011100100000"; -- -0.068577341735363
	pesos_i(9358) := b"1111111111111111_1111111111111111_1100110110111011_1110101101000000"; -- -0.1963513344526291
	pesos_i(9359) := b"0000000000000000_0000000000000000_0000110010001111_0010011011000000"; -- 0.049059316515922546
	pesos_i(9360) := b"0000000000000000_0000000000000000_0101010011001001_0001011110000000"; -- 0.3311934173107147
	pesos_i(9361) := b"1111111111111111_1111111111111111_1101101111110010_0100001011000000"; -- -0.14083464443683624
	pesos_i(9362) := b"1111111111111111_1111111111111111_1001011110110001_1010010110000000"; -- -0.4074455797672272
	pesos_i(9363) := b"1111111111111111_1111111111111111_1010100001001110_0001011010000000"; -- -0.34255847334861755
	pesos_i(9364) := b"0000000000000000_0000000000000000_0000001001001010_1010001001010000"; -- 0.008951324969530106
	pesos_i(9365) := b"1111111111111111_1111111111111111_1010110110001000_0111111010000000"; -- -0.3221360146999359
	pesos_i(9366) := b"1111111111111111_1111111111111111_1110110100100011_1011100000100000"; -- -0.07367371767759323
	pesos_i(9367) := b"1111111111111111_1111111111111111_1111010111100100_1101011001110000"; -- -0.03947696462273598
	pesos_i(9368) := b"0000000000000000_0000000000000000_0101000111001000_1010000010000000"; -- 0.31946757435798645
	pesos_i(9369) := b"1111111111111111_1111111111111111_1100101110010110_0001100111000000"; -- -0.20474089682102203
	pesos_i(9370) := b"1111111111111111_1111111111111111_1011000101101101_1010001110000000"; -- -0.3069207966327667
	pesos_i(9371) := b"0000000000000000_0000000000000000_0111011011110010_0110101010000000"; -- 0.4646364748477936
	pesos_i(9372) := b"0000000000000000_0000000000000000_0000000111110001_0111000110010110"; -- 0.007590388413518667
	pesos_i(9373) := b"1111111111111111_1111111111111111_1010110111001100_0100001110000000"; -- -0.32110193371772766
	pesos_i(9374) := b"0000000000000000_0000000000000000_0110100100110110_1111101100000000"; -- 0.4109951853752136
	pesos_i(9375) := b"1111111111111111_1111111111111111_1101000111111001_0100001111000000"; -- -0.17979027330875397
	pesos_i(9376) := b"0000000000000000_0000000000000000_0111000111100011_1111110010000000"; -- 0.4448850452899933
	pesos_i(9377) := b"1111111111111111_1111111111111111_1011000010011000_1011110000000000"; -- -0.3101694583892822
	pesos_i(9378) := b"1111111111111111_1111111111111111_1111110011100100_0000101111100000"; -- -0.012145288288593292
	pesos_i(9379) := b"0000000000000000_0000000000000000_0010011110011000_1110101011000000"; -- 0.15467707812786102
	pesos_i(9380) := b"1111111111111111_1111111111111111_0010010100001001_1010010000000000"; -- -0.8553216457366943
	pesos_i(9381) := b"0000000000000000_0000000000000000_0111001000101001_1100001010000000"; -- 0.4459497034549713
	pesos_i(9382) := b"1111111111111111_1111111111111111_0110001100100111_0000011000000000"; -- -0.6126857995986938
	pesos_i(9383) := b"0000000000000000_0000000000000000_0100111100000000_0001100110000000"; -- 0.3085952699184418
	pesos_i(9384) := b"0000000000000000_0000000000000000_0010000111111101_1001001111000000"; -- 0.13277553021907806
	pesos_i(9385) := b"0000000000000000_0000000000000000_0111101000111110_0111011100000000"; -- 0.47751563787460327
	pesos_i(9386) := b"1111111111111111_1111111111111111_1111010100010111_1010001100110000"; -- -0.042608071118593216
	pesos_i(9387) := b"1111111111111111_1111111111111111_1110111100101101_1110011001000000"; -- -0.06570588052272797
	pesos_i(9388) := b"1111111111111111_1111111111111111_0001000110000010_0010101100000000"; -- -0.9316075444221497
	pesos_i(9389) := b"1111111111111111_1111111111111111_1111111001011111_1000010000010110"; -- -0.006355042103677988
	pesos_i(9390) := b"1111111111111111_1111111111111111_1110000100001100_1010111000100000"; -- -0.12090026587247849
	pesos_i(9391) := b"1111111111111111_1111111111111111_1111000110011001_1111000111110000"; -- -0.056244734674692154
	pesos_i(9392) := b"0000000000000000_0000000000000000_0010000110111000_0000001011000000"; -- 0.13171403110027313
	pesos_i(9393) := b"0000000000000000_0000000000000000_0000111111001101_0110001110000000"; -- 0.06172773241996765
	pesos_i(9394) := b"0000000000000000_0000000000000000_0011101110100001_0100010001000000"; -- 0.23292948305606842
	pesos_i(9395) := b"0000000000000000_0000000000000000_0000001011101010_1110011110101100"; -- 0.011396865360438824
	pesos_i(9396) := b"0000000000000000_0000000000000000_0100100100001000_0101110100000000"; -- 0.2852838635444641
	pesos_i(9397) := b"1111111111111111_1111111111111111_1001111111001111_0010011010000000"; -- -0.37574538588523865
	pesos_i(9398) := b"0000000000000000_0000000000000000_0101100011110101_0011110100000000"; -- 0.3474920392036438
	pesos_i(9399) := b"1111111111111111_1111111111111111_1001100101010011_0000100100000000"; -- -0.4010767340660095
	pesos_i(9400) := b"1111111111111111_1111111111111111_1010010100001001_0011011010000000"; -- -0.35532817244529724
	pesos_i(9401) := b"1111111111111111_1111111111111111_1010000001000100_0000000000000000"; -- -0.37396240234375
	pesos_i(9402) := b"0000000000000000_0000000000000000_0011110111110110_1101010111000000"; -- 0.24204765260219574
	pesos_i(9403) := b"1111111111111111_1111111111111111_1101110011010100_1001000111000000"; -- -0.137381449341774
	pesos_i(9404) := b"0000000000000000_0000000000000000_0001000100101110_1100111000000000"; -- 0.06712043285369873
	pesos_i(9405) := b"0000000000000000_0000000000000000_0101010101010111_0001000100000000"; -- 0.3333597779273987
	pesos_i(9406) := b"1111111111111111_1111111111111111_1010010001110111_0001001110000000"; -- -0.3575580418109894
	pesos_i(9407) := b"1111111111111111_1111111111111111_1101000000111111_1001010101000000"; -- -0.18652980029582977
	pesos_i(9408) := b"0000000000000000_0000000000000000_0000111100001110_1111100011000000"; -- 0.05882219970226288
	pesos_i(9409) := b"0000000000000000_0000000000000000_0011011111010111_1011100010000000"; -- 0.21813538670539856
	pesos_i(9410) := b"1111111111111111_1111111111111111_0111101111011011_0100111100000000"; -- -0.5161848664283752
	pesos_i(9411) := b"1111111111111111_1111111111111111_1010111011100001_1110100100000000"; -- -0.31686538457870483
	pesos_i(9412) := b"1111111111111111_1111111111111111_1110111110001100_1101111100100000"; -- -0.06425672024488449
	pesos_i(9413) := b"0000000000000000_0000000000000000_0011011101001110_1101110011000000"; -- 0.21604709327220917
	pesos_i(9414) := b"1111111111111111_1111111111111111_1011110001001101_0011010010000000"; -- -0.2644469439983368
	pesos_i(9415) := b"1111111111111111_1111111111111111_1010001011011010_1001001100000000"; -- -0.363852322101593
	pesos_i(9416) := b"0000000000000000_0000000000000000_0001110001001100_1011011011100000"; -- 0.1105455681681633
	pesos_i(9417) := b"1111111111111111_1111111111111111_1100100000110100_0010011011000000"; -- -0.21795423328876495
	pesos_i(9418) := b"0000000000000000_0000000000000000_0100100101100011_0111101110000000"; -- 0.28667423129081726
	pesos_i(9419) := b"1111111111111111_1111111111111111_1000110001000011_1010010100000000"; -- -0.45209282636642456
	pesos_i(9420) := b"1111111111111111_1111111111111111_1111100001000100_0010010110100000"; -- -0.030210159718990326
	pesos_i(9421) := b"0000000000000000_0000000000000000_0001110100011001_0000000011100000"; -- 0.11366277188062668
	pesos_i(9422) := b"1111111111111111_1111111111111111_1011111101011011_1101000100000000"; -- -0.25250524282455444
	pesos_i(9423) := b"1111111111111111_1111111111111111_1110101100110101_0101101011000000"; -- -0.08121712505817413
	pesos_i(9424) := b"1111111111111111_1111111111111111_0111001000111001_1010010100000000"; -- -0.5538079142570496
	pesos_i(9425) := b"0000000000000000_0000000000000000_0001001011111100_0111000010100000"; -- 0.07416442781686783
	pesos_i(9426) := b"0000000000000000_0000000000000000_0011111110111011_1100101011000000"; -- 0.2489592283964157
	pesos_i(9427) := b"1111111111111111_1111111111111111_1101001010100011_1000110101000000"; -- -0.17719189822673798
	pesos_i(9428) := b"1111111111111111_1111111111111111_1011010001000100_0001111010000000"; -- -0.29583558440208435
	pesos_i(9429) := b"0000000000000000_0000000000000000_0010001101101001_1010010010000000"; -- 0.13833072781562805
	pesos_i(9430) := b"1111111111111111_1111111111111111_1101000001011000_1010011000000000"; -- -0.18614733219146729
	pesos_i(9431) := b"0000000000000000_0000000000000000_0100010101001101_0011100000000000"; -- 0.2707095146179199
	pesos_i(9432) := b"0000000000000000_0000000000000000_0110010101101011_0111101110000000"; -- 0.39617130160331726
	pesos_i(9433) := b"0000000000000000_0000000000000000_1000010000001100_0000110100000000"; -- 0.5158088803291321
	pesos_i(9434) := b"1111111111111111_1111111111111111_0110000100011001_1101110100000000"; -- -0.6206991076469421
	pesos_i(9435) := b"1111111111111111_1111111111111111_1011010100111001_1011010010000000"; -- -0.29208824038505554
	pesos_i(9436) := b"1111111111111111_1111111111111111_1101011010101110_1111010110000000"; -- -0.16139283776283264
	pesos_i(9437) := b"0000000000000000_0000000000000000_0011011001110001_0000100011000000"; -- 0.21266226470470428
	pesos_i(9438) := b"0000000000000000_0000000000000000_0110100100001111_1000000110000000"; -- 0.4103928506374359
	pesos_i(9439) := b"0000000000000000_0000000000000000_0000100011001001_1001110100000000"; -- 0.034326374530792236
	pesos_i(9440) := b"1111111111111111_1111111111111111_1001000101100011_1100100000000000"; -- -0.4320712089538574
	pesos_i(9441) := b"1111111111111111_1111111111111111_0100011100000011_1101110000000000"; -- -0.7225973606109619
	pesos_i(9442) := b"0000000000000000_0000000000000000_0010000101001001_1111101000000000"; -- 0.13003504276275635
	pesos_i(9443) := b"0000000000000000_0000000000000000_0011000001110111_1100001111000000"; -- 0.18932746350765228
	pesos_i(9444) := b"1111111111111111_1111111111111111_1011100001000101_1100011100000000"; -- -0.2801852822303772
	pesos_i(9445) := b"1111111111111111_1111111111111111_1111111010110011_0110000110111110"; -- -0.005075350869446993
	pesos_i(9446) := b"0000000000000000_0000000000000000_0010011011110101_1100011111000000"; -- 0.15218780934810638
	pesos_i(9447) := b"1111111111111111_1111111111111111_0111101011010001_1110000100000000"; -- -0.520235002040863
	pesos_i(9448) := b"1111111111111111_1111111111111111_1110011001100000_0100000100100000"; -- -0.100093774497509
	pesos_i(9449) := b"1111111111111111_1111111111111111_1101111001110000_0011010100000000"; -- -0.1311003565788269
	pesos_i(9450) := b"1111111111111111_1111111111111111_1110111000010011_1100110001100000"; -- -0.07001040130853653
	pesos_i(9451) := b"0000000000000000_0000000000000000_0100100101001110_1101000110000000"; -- 0.28635892271995544
	pesos_i(9452) := b"1111111111111111_1111111111111111_0010001110110110_0101110100000000"; -- -0.8604986071586609
	pesos_i(9453) := b"1111111111111111_1111111111111111_1101001111111010_0110110010000000"; -- -0.17196008563041687
	pesos_i(9454) := b"1111111111111111_1111111111111111_1110110101000000_0101111100000000"; -- -0.07323652505874634
	pesos_i(9455) := b"0000000000000000_0000000000000000_1001011111010111_0100110000000000"; -- 0.5931289196014404
	pesos_i(9456) := b"0000000000000000_0000000000000000_0011110011011011_0001000110000000"; -- 0.23771771788597107
	pesos_i(9457) := b"0000000000000000_0000000000000000_0110011101000011_1011111100000000"; -- 0.4033774733543396
	pesos_i(9458) := b"1111111111111111_1111111111111111_0110111100111110_0010001100000000"; -- -0.5654581189155579
	pesos_i(9459) := b"1111111111111111_1111111111111110_1111100000101010_1001000000000000"; -- -1.0306005477905273
	pesos_i(9460) := b"0000000000000000_0000000000000000_0000011010010101_1000001111001000"; -- 0.025718914344906807
	pesos_i(9461) := b"0000000000000000_0000000000000000_0110100111100110_1010000100000000"; -- 0.41367536783218384
	pesos_i(9462) := b"0000000000000000_0000000000000000_0000110111111010_0011111101100000"; -- 0.05459972470998764
	pesos_i(9463) := b"1111111111111111_1111111111111111_1100010011000111_1111100110000000"; -- -0.23132362961769104
	pesos_i(9464) := b"0000000000000000_0000000000000000_0011011101010110_0000011011000000"; -- 0.21615640819072723
	pesos_i(9465) := b"0000000000000000_0000000000000000_0000011100011011_1010111100111000"; -- 0.027766181156039238
	pesos_i(9466) := b"1111111111111111_1111111111111111_0101100101010011_0010111000000000"; -- -0.6510745286941528
	pesos_i(9467) := b"1111111111111111_1111111111111111_1011101101010101_1110101010000000"; -- -0.26822027564048767
	pesos_i(9468) := b"1111111111111111_1111111111111111_0110010110110001_0100111000000000"; -- -0.602763295173645
	pesos_i(9469) := b"0000000000000000_0000000000000000_0010010010100011_0000110001000000"; -- 0.143112912774086
	pesos_i(9470) := b"1111111111111111_1111111111111111_1100101001111101_1111101100000000"; -- -0.20901519060134888
	pesos_i(9471) := b"0000000000000000_0000000000000000_0100110111111101_0100100000000000"; -- 0.30464601516723633

    return pesos_i;
    end function;
end package body mnist_weights;
    