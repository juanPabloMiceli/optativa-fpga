
-- ARCHIVO AUTOGENERADO CON model/tensorflow_model.py

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.perceptron_package.perceptron_input;

package mnist_inputs_9 is
    function GetInputs(Dummy: natural)
    return perceptron_input;
end package mnist_inputs_9;

package body mnist_inputs_9 is
    function GetInputs(Dummy: natural) return perceptron_input is
        variable pesos_i : perceptron_input(63 downto 0);
    begin
	pesos_i(0) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(1) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(2) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(3) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(4) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(5) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(6) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(7) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(8) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(9) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(10) := b"0000000000000000_0000000000000000_0011010010010010_1100011010101101"; -- 0.20536462529984795
	pesos_i(11) := b"0000000000000000_0000000000000000_0111101110100100_0000000000011011"; -- 0.48297119777026437
	pesos_i(12) := b"0000000000000000_0000000000000000_0000011010011111_0010101011110110"; -- 0.025866208084564236
	pesos_i(13) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(14) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(15) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(16) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(17) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(18) := b"0000000000000000_0000000000000000_1101110000100110_1001111111110110"; -- 0.8599643684431133
	pesos_i(19) := b"0000000000000000_0000000000000000_0111101010100110_1100100011001111"; -- 0.47910742818810226
	pesos_i(20) := b"0000000000000000_0000000000000000_0101111010011000_1010111011011100"; -- 0.36951725835091764
	pesos_i(21) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(22) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(23) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(24) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(25) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(26) := b"0000000000000000_0000000000000000_0111001100000001_0001001010011011"; -- 0.4492351178434174
	pesos_i(27) := b"0000000000000000_0000000000000000_1000101001111010_0011110110001111"; -- 0.5409277415026961
	pesos_i(28) := b"0000000000000000_0000000000000000_1000100000111000_0000011000001001"; -- 0.5321048520253214
	pesos_i(29) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(30) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(31) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(32) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(33) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(34) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(35) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(36) := b"0000000000000000_0000000000000000_0110010100110111_1101100111010010"; -- 0.3953834664354819
	pesos_i(37) := b"0000000000000000_0000000000000000_0100011010010110_0100111011011000"; -- 0.27573101772605496
	pesos_i(38) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(39) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(40) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(41) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(42) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(43) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(44) := b"0000000000000000_0000000000000000_0100011011110010_1000001100100101"; -- 0.27713794376318823
	pesos_i(45) := b"0000000000000000_0000000000000000_1011101100110101_1001100101110100"; -- 0.7312866122299719
	pesos_i(46) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(47) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(48) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(49) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(50) := b"0000000000000000_0000000000000000_0010000011011011_1011110000101100"; -- 0.12835289081240497
	pesos_i(51) := b"0000000000000000_0000000000000000_0111111010011011_1010010111111111"; -- 0.4945625065167507
	pesos_i(52) := b"0000000000000000_0000000000000000_1001010010000100_0011000101000000"; -- 0.5801420956109407
	pesos_i(53) := b"0000000000000000_0000000000000000_1001111110010110_1001101111111110"; -- 0.6233918661632547
	pesos_i(54) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(55) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(56) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(57) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(58) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(59) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(60) := b"0000000000000000_0000000000000000_0001100110001010_1000000100100010"; -- 0.09976965975474776
	pesos_i(61) := b"0000000000000000_0000000000000000_0000011000100011_0101010011000101"; -- 0.02397661023704826
	pesos_i(62) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0
	pesos_i(63) := b"0000000000000000_0000000000000000_0000000000000000_0000000000000000"; -- 0.0

    return pesos_i;
    end function;
end package body mnist_inputs_9;
    